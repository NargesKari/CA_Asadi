/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
alop
**
**
**
*****************************************************************************/
module
alop(
func,
oooo,
op
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[5:0]
func;
input
[5:0]
op;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[3:0]
oooo;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[3:0]
s_logisimBus11;
wire
[5:0]
s_logisimBus15;
wire
[5:0]
s_logisimBus17;
wire
[5:0]
s_logisimBus29;
wire
[5:0]
s_logisimBus35;
wire
[5:0]
s_logisimBus36;
wire
[5:0]
s_logisimBus39;
wire
[5:0]
s_logisimBus43;
wire
[5:0]
s_logisimBus47;
wire
[5:0]
s_logisimBus5;
wire
[5:0]
s_logisimBus53;
wire
[5:0]
s_logisimBus55;
wire
[5:0]
s_logisimBus57;
wire
[5:0]
s_logisimBus61;
wire
[5:0]
s_logisimBus65;
wire
[5:0]
s_logisimBus68;
wire
[5:0]
s_logisimBus73;
wire
[5:0]
s_logisimBus76;
wire
[5:0]
s_logisimBus83;
wire
[5:0]
s_logisimBus9;
wire
[5:0]
s_logisimBus91;
wire
[5:0]
s_logisimBus92;
wire
[5:0]
s_logisimBus94;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet10;
wire
s_logisimNet12;
wire
s_logisimNet13;
wire
s_logisimNet14;
wire
s_logisimNet16;
wire
s_logisimNet18;
wire
s_logisimNet19;
wire
s_logisimNet2;
wire
s_logisimNet20;
wire
s_logisimNet21;
wire
s_logisimNet22;
wire
s_logisimNet23;
wire
s_logisimNet24;
wire
s_logisimNet25;
wire
s_logisimNet26;
wire
s_logisimNet27;
wire
s_logisimNet28;
wire
s_logisimNet3;
wire
s_logisimNet30;
wire
s_logisimNet31;
wire
s_logisimNet32;
wire
s_logisimNet33;
wire
s_logisimNet34;
wire
s_logisimNet37;
wire
s_logisimNet38;
wire
s_logisimNet4;
wire
s_logisimNet40;
wire
s_logisimNet41;
wire
s_logisimNet42;
wire
s_logisimNet44;
wire
s_logisimNet45;
wire
s_logisimNet46;
wire
s_logisimNet48;
wire
s_logisimNet49;
wire
s_logisimNet50;
wire
s_logisimNet51;
wire
s_logisimNet52;
wire
s_logisimNet54;
wire
s_logisimNet56;
wire
s_logisimNet58;
wire
s_logisimNet59;
wire
s_logisimNet6;
wire
s_logisimNet60;
wire
s_logisimNet62;
wire
s_logisimNet63;
wire
s_logisimNet64;
wire
s_logisimNet66;
wire
s_logisimNet67;
wire
s_logisimNet69;
wire
s_logisimNet7;
wire
s_logisimNet70;
wire
s_logisimNet71;
wire
s_logisimNet72;
wire
s_logisimNet74;
wire
s_logisimNet75;
wire
s_logisimNet77;
wire
s_logisimNet78;
wire
s_logisimNet79;
wire
s_logisimNet8;
wire
s_logisimNet80;
wire
s_logisimNet81;
wire
s_logisimNet82;
wire
s_logisimNet84;
wire
s_logisimNet85;
wire
s_logisimNet86;
wire
s_logisimNet87;
wire
s_logisimNet88;
wire
s_logisimNet89;
wire
s_logisimNet90;
wire
s_logisimNet93;
wire
s_logisimNet95;
wire
s_logisimNet96;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus55[5:0]
=
op;
assign
s_logisimBus9[5:0]
=
func;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
oooo
=
s_logisimBus11[3:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus5[5:0]
=
{2'b10,
4'h2};
assign
s_logisimBus65[5:0]
=
{2'b10,
4'h0};
assign
s_logisimBus43[5:0]
=
{2'b10,
4'h0};
assign
s_logisimBus57[5:0]
=
{2'b10,
4'h4};
assign
s_logisimBus29[5:0]
=
{2'b10,
4'h2};
assign
s_logisimBus76[5:0]
=
{2'b10,
4'h0};
assign
s_logisimBus47[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus53[5:0]
=
{2'b10,
4'h5};
assign
s_logisimBus91[5:0]
=
{2'b00,
4'h6};
assign
s_logisimBus94[5:0]
=
{2'b10,
4'h5};
assign
s_logisimBus73[5:0]
=
{2'b10,
4'h4};
assign
s_logisimBus35[5:0]
=
{2'b00,
4'h6};
assign
s_logisimBus15[5:0]
=
{2'b00,
4'h4};
assign
s_logisimBus61[5:0]
=
{2'b10,
4'h6};
assign
s_logisimBus36[5:0]
=
{2'b10,
4'h4};
assign
s_logisimBus68[5:0]
=
{2'b10,
4'h2};
assign
s_logisimBus39[5:0]
=
{2'b10,
4'h6};
assign
s_logisimNet26
=
1'b1;
assign
s_logisimNet32
=
1'b0;
assign
s_logisimBus83[5:0]
=
{2'b00,
4'h7};
assign
s_logisimNet80
=
1'b1;
assign
s_logisimNet22
=
1'b0;
assign
s_logisimBus17[5:0]
=
{2'b10,
4'h0};
assign
s_logisimBus92[5:0]
=
{2'b00,
4'h4};
assign
s_logisimNet48
=
1'b1;
assign
s_logisimNet52
=
1'b0;
assign
s_logisimNet89
=
1'b1;
assign
s_logisimNet1
=
1'b0;
assign
s_logisimNet46
=
~s_logisimNet74;
assign
s_logisimNet37
=
~s_logisimNet74;
assign
s_logisimNet23
=
~s_logisimNet74;
assign
s_logisimNet2
=
~s_logisimNet74;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE
#(.BubblesMask(2'b00))
GATES_1
(.input1(s_logisimNet93),
.input2(s_logisimNet90),
.result(s_logisimNet8));
AND_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet74),
.input2(s_logisimNet19),
.result(s_logisimNet58));
AND_GATE
#(.BubblesMask(2'b00))
GATES_3
(.input1(s_logisimNet74),
.input2(s_logisimNet20),
.result(s_logisimNet45));
AND_GATE
#(.BubblesMask(2'b00))
GATES_4
(.input1(s_logisimNet74),
.input2(s_logisimNet77),
.result(s_logisimNet54));
AND_GATE
#(.BubblesMask(2'b00))
GATES_5
(.input1(s_logisimNet74),
.input2(s_logisimNet78),
.result(s_logisimNet87));
AND_GATE
#(.BubblesMask(2'b00))
GATES_6
(.input1(s_logisimNet74),
.input2(s_logisimNet95),
.result(s_logisimNet50));
AND_GATE
#(.BubblesMask(2'b00))
GATES_7
(.input1(s_logisimNet74),
.input2(s_logisimNet96),
.result(s_logisimNet24));
AND_GATE
#(.BubblesMask(2'b00))
GATES_8
(.input1(s_logisimNet74),
.input2(s_logisimNet84),
.result(s_logisimNet6));
AND_GATE
#(.BubblesMask(2'b00))
GATES_9
(.input1(s_logisimNet74),
.input2(s_logisimNet85),
.result(s_logisimNet4));
AND_GATE
#(.BubblesMask(2'b00))
GATES_10
(.input1(s_logisimNet74),
.input2(s_logisimNet66),
.result(s_logisimNet69));
AND_GATE
#(.BubblesMask(2'b00))
GATES_11
(.input1(s_logisimNet74),
.input2(s_logisimNet3),
.result(s_logisimNet7));
OR_GATE
#(.BubblesMask(2'b00))
GATES_12
(.input1(s_logisimNet58),
.input2(s_logisimNet45),
.result(s_logisimNet25));
AND_GATE
#(.BubblesMask(2'b00))
GATES_13
(.input1(s_logisimNet74),
.input2(s_logisimNet28),
.result(s_logisimNet33));
AND_GATE
#(.BubblesMask(2'b00))
GATES_14
(.input1(s_logisimNet74),
.input2(s_logisimNet10),
.result(s_logisimNet75));
AND_GATE
#(.BubblesMask(2'b00))
GATES_15
(.input1(s_logisimNet74),
.input2(s_logisimNet56),
.result(s_logisimNet59));
OR_GATE
#(.BubblesMask(2'b00))
GATES_16
(.input1(s_logisimNet54),
.input2(s_logisimNet87),
.result(s_logisimNet63));
AND_GATE
#(.BubblesMask(2'b00))
GATES_17
(.input1(s_logisimNet74),
.input2(s_logisimNet30),
.result(s_logisimNet16));
OR_GATE
#(.BubblesMask(2'b00))
GATES_18
(.input1(s_logisimNet25),
.input2(s_logisimNet75),
.result(s_logisimNet71));
OR_GATE
#(.BubblesMask(2'b00))
GATES_19
(.input1(s_logisimNet50),
.input2(s_logisimNet24),
.result(s_logisimNet0));
OR_GATE
#(.BubblesMask(2'b00))
GATES_20
(.input1(s_logisimNet6),
.input2(s_logisimNet4),
.result(s_logisimNet72));
AND_GATE
#(.BubblesMask(2'b00))
GATES_21
(.input1(s_logisimNet74),
.input2(s_logisimNet67),
.result(s_logisimNet64));
AND_GATE
#(.BubblesMask(2'b00))
GATES_22
(.input1(s_logisimNet74),
.input2(s_logisimNet51),
.result(s_logisimNet41));
OR_GATE
#(.BubblesMask(2'b00))
GATES_23
(.input1(s_logisimNet63),
.input2(s_logisimNet16),
.result(s_logisimNet14));
OR_GATE
#(.BubblesMask(2'b00))
GATES_24
(.input1(s_logisimNet71),
.input2(s_logisimNet69),
.result(s_logisimNet21));
OR_GATE
#(.BubblesMask(2'b00))
GATES_25
(.input1(s_logisimNet0),
.input2(s_logisimNet64),
.result(s_logisimNet62));
OR_GATE
#(.BubblesMask(2'b00))
GATES_26
(.input1(s_logisimNet72),
.input2(s_logisimNet41),
.result(s_logisimNet40));
OR_GATE
#(.BubblesMask(2'b00))
GATES_27
(.input1(s_logisimNet14),
.input2(s_logisimNet7),
.result(s_logisimNet79));
OR_GATE
#(.BubblesMask(2'b00))
GATES_28
(.input1(s_logisimNet21),
.input2(s_logisimNet46),
.result(s_logisimNet44));
OR_GATE
#(.BubblesMask(2'b00))
GATES_29
(.input1(s_logisimNet62),
.input2(s_logisimNet59),
.result(s_logisimNet34));
OR_GATE
#(.BubblesMask(2'b00))
GATES_30
(.input1(s_logisimNet40),
.input2(s_logisimNet33),
.result(s_logisimNet88));
OR_GATE
#(.BubblesMask(2'b00))
GATES_31
(.input1(s_logisimNet79),
.input2(s_logisimNet37),
.result(s_logisimNet86));
AND_GATE
#(.BubblesMask(2'b00))
GATES_32
(.input1(s_logisimNet74),
.input2(s_logisimNet13),
.result(s_logisimNet31));
OR_GATE
#(.BubblesMask(2'b00))
GATES_33
(.input1(s_logisimNet34),
.input2(s_logisimNet23),
.result(s_logisimNet12));
OR_GATE
#(.BubblesMask(2'b00))
GATES_34
(.input1(s_logisimNet88),
.input2(s_logisimNet2),
.result(s_logisimNet93));
AND_GATE
#(.BubblesMask(2'b00))
GATES_35
(.input1(s_logisimNet74),
.input2(s_logisimNet70),
.result(s_logisimNet81));
OR_GATE
#(.BubblesMask(2'b00))
GATES_36
(.input1(s_logisimNet44),
.input2(s_logisimNet31),
.result(s_logisimNet42));
AND_GATE
#(.BubblesMask(2'b00))
GATES_37
(.input1(s_logisimNet74),
.input2(s_logisimNet82),
.result(s_logisimNet90));
OR_GATE
#(.BubblesMask(2'b00))
GATES_38
(.input1(s_logisimNet86),
.input2(s_logisimNet81),
.result(s_logisimNet27));
Multiplexer_2
PLEXERS_39
(.enable(1'b1),
.muxIn_0(s_logisimNet26),
.muxIn_1(s_logisimNet32),
.muxOut(s_logisimBus11[3]),
.sel(s_logisimNet42));
Multiplexer_2
PLEXERS_40
(.enable(1'b1),
.muxIn_0(s_logisimNet80),
.muxIn_1(s_logisimNet22),
.muxOut(s_logisimBus11[2]),
.sel(s_logisimNet27));
Multiplexer_2
PLEXERS_41
(.enable(1'b1),
.muxIn_0(s_logisimNet48),
.muxIn_1(s_logisimNet52),
.muxOut(s_logisimBus11[0]),
.sel(s_logisimNet12));
Multiplexer_2
PLEXERS_42
(.enable(1'b1),
.muxIn_0(s_logisimNet89),
.muxIn_1(s_logisimNet1),
.muxOut(s_logisimBus11[1]),
.sel(s_logisimNet8));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_43
(.aEqualsB(s_logisimNet19),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus76[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_44
(.aEqualsB(s_logisimNet20),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus68[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_45
(.aEqualsB(s_logisimNet77),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus17[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_46
(.aEqualsB(s_logisimNet78),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus5[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_47
(.aEqualsB(s_logisimNet95),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus65[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_48
(.aEqualsB(s_logisimNet96),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus57[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_49
(.aEqualsB(s_logisimNet84),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus43[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_50
(.aEqualsB(s_logisimNet85),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus29[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_51
(.aEqualsB(s_logisimNet66),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus53[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_52
(.aEqualsB(s_logisimNet74),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus55[5:0]),
.dataB(s_logisimBus47[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_53
(.aEqualsB(s_logisimNet3),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus91[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_54
(.aEqualsB(s_logisimNet10),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus73[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_55
(.aEqualsB(s_logisimNet28),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus94[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_56
(.aEqualsB(s_logisimNet56),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus35[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_57
(.aEqualsB(s_logisimNet30),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_58
(.aEqualsB(s_logisimNet67),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus61[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_59
(.aEqualsB(s_logisimNet51),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus36[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_60
(.aEqualsB(s_logisimNet13),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus39[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_61
(.aEqualsB(s_logisimNet70),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus83[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(1))
ARITH_62
(.aEqualsB(s_logisimNet82),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus92[5:0]));
endmodule