/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
PC_Update
**
**
**
*****************************************************************************/
module
PC_Update(
Branch,
Eq,
Imm,
Jump,
PC,
PC_out,
divIsActive,
isNe
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
Branch;
input
[31:0]
Eq;
input
[15:0]
Imm;
input
Jump;
input
[8:0]
PC;
input
divIsActive;
input
isNe;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[8:0]
PC_out;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[15:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus11;
wire
[8:0]
s_logisimBus13;
wire
[8:0]
s_logisimBus14;
wire
[8:0]
s_logisimBus16;
wire
[31:0]
s_logisimBus19;
wire
[8:0]
s_logisimBus2;
wire
[8:0]
s_logisimBus4;
wire
[8:0]
s_logisimBus5;
wire
[8:0]
s_logisimBus8;
wire
s_logisimNet10;
wire
s_logisimNet12;
wire
s_logisimNet15;
wire
s_logisimNet17;
wire
s_logisimNet18;
wire
s_logisimNet3;
wire
s_logisimNet6;
wire
s_logisimNet7;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus0[15:0]
=
Imm;
assign
s_logisimBus11[31:0]
=
Eq;
assign
s_logisimBus2[8:0]
=
PC;
assign
s_logisimNet10
=
isNe;
assign
s_logisimNet3
=
divIsActive;
assign
s_logisimNet6
=
Branch;
assign
s_logisimNet7
=
Jump;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
PC_out
=
s_logisimBus16[8:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus14[8:0]
=
{1'b0,
8'h01};
assign
s_logisimNet17
=
1'b0;
assign
s_logisimBus19[31:0]
=
32'h00000000;
assign
s_logisimNet18
=
1'b0;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
XOR_GATE_ONEHOT
#(.BubblesMask(2'b00))
GATES_1
(.input1(s_logisimNet10),
.input2(s_logisimNet9),
.result(s_logisimNet15));
AND_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet6),
.input2(s_logisimNet15),
.result(s_logisimNet12));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus5[8:0]),
.muxIn_1(s_logisimBus8[8:0]),
.muxOut(s_logisimBus4[8:0]),
.sel(s_logisimNet12));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus4[8:0]),
.muxIn_1(s_logisimBus0[8:0]),
.muxOut(s_logisimBus13[8:0]),
.sel(s_logisimNet7));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus13[8:0]),
.muxIn_1(s_logisimBus2[8:0]),
.muxOut(s_logisimBus16[8:0]),
.sel(s_logisimNet3));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_6
(.carryIn(s_logisimNet17),
.carryOut(),
.dataA(s_logisimBus14[8:0]),
.dataB(s_logisimBus2[8:0]),
.result(s_logisimBus5[8:0]));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_7
(.carryIn(s_logisimNet18),
.carryOut(),
.dataA(s_logisimBus5[8:0]),
.dataB(s_logisimBus0[8:0]),
.result(s_logisimBus8[8:0]));
Comparator
#(.nrOfBits(32),
.twosComplement(1))
ARITH_8
(.aEqualsB(s_logisimNet9),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus11[31:0]),
.dataB(s_logisimBus19[31:0]));
endmodule