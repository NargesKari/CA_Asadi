/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
divi
**
**
**
*****************************************************************************/
module
divi(
clk,
dividend,
divisor,
done,
quotient,
remainder
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
clk;
input
[31:0]
dividend;
input
[31:0]
divisor;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
done;
output
[31:0]
quotient;
output
[31:0]
remainder;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[63:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus1;
wire
[31:0]
s_logisimBus10;
wire
[31:0]
s_logisimBus13;
wire
[31:0]
s_logisimBus18;
wire
[31:0]
s_logisimBus19;
wire
[31:0]
s_logisimBus20;
wire
[31:0]
s_logisimBus21;
wire
[63:0]
s_logisimBus25;
wire
[31:0]
s_logisimBus27;
wire
[63:0]
s_logisimBus28;
wire
[63:0]
s_logisimBus29;
wire
[31:0]
s_logisimBus3;
wire
[31:0]
s_logisimBus32;
wire
[30:0]
s_logisimBus34;
wire
[63:0]
s_logisimBus35;
wire
[31:0]
s_logisimBus36;
wire
[31:0]
s_logisimBus4;
wire
[63:0]
s_logisimBus5;
wire
[31:0]
s_logisimBus6;
wire
[30:0]
s_logisimBus9;
wire
s_logisimNet11;
wire
s_logisimNet12;
wire
s_logisimNet14;
wire
s_logisimNet15;
wire
s_logisimNet16;
wire
s_logisimNet17;
wire
s_logisimNet2;
wire
s_logisimNet22;
wire
s_logisimNet23;
wire
s_logisimNet24;
wire
s_logisimNet26;
wire
s_logisimNet30;
wire
s_logisimNet31;
wire
s_logisimNet33;
wire
s_logisimNet37;
wire
s_logisimNet38;
wire
s_logisimNet39;
wire
s_logisimNet7;
wire
s_logisimNet8;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
wiring
is
defined
**
*******************************************************************************/
assign
s_logisimBus21[10]
=
s_logisimBus9[9];
assign
s_logisimBus21[11]
=
s_logisimBus9[10];
assign
s_logisimBus21[12]
=
s_logisimBus9[11];
assign
s_logisimBus21[13]
=
s_logisimBus9[12];
assign
s_logisimBus21[14]
=
s_logisimBus9[13];
assign
s_logisimBus21[15]
=
s_logisimBus9[14];
assign
s_logisimBus21[16]
=
s_logisimBus9[15];
assign
s_logisimBus21[17]
=
s_logisimBus9[16];
assign
s_logisimBus21[18]
=
s_logisimBus9[17];
assign
s_logisimBus21[19]
=
s_logisimBus9[18];
assign
s_logisimBus21[1]
=
s_logisimBus9[0];
assign
s_logisimBus21[20]
=
s_logisimBus9[19];
assign
s_logisimBus21[21]
=
s_logisimBus9[20];
assign
s_logisimBus21[22]
=
s_logisimBus9[21];
assign
s_logisimBus21[23]
=
s_logisimBus9[22];
assign
s_logisimBus21[24]
=
s_logisimBus9[23];
assign
s_logisimBus21[25]
=
s_logisimBus9[24];
assign
s_logisimBus21[26]
=
s_logisimBus9[25];
assign
s_logisimBus21[27]
=
s_logisimBus9[26];
assign
s_logisimBus21[28]
=
s_logisimBus9[27];
assign
s_logisimBus21[29]
=
s_logisimBus9[28];
assign
s_logisimBus21[2]
=
s_logisimBus9[1];
assign
s_logisimBus21[30]
=
s_logisimBus9[29];
assign
s_logisimBus21[31]
=
s_logisimBus9[30];
assign
s_logisimBus21[3]
=
s_logisimBus9[2];
assign
s_logisimBus21[4]
=
s_logisimBus9[3];
assign
s_logisimBus21[5]
=
s_logisimBus9[4];
assign
s_logisimBus21[6]
=
s_logisimBus9[5];
assign
s_logisimBus21[7]
=
s_logisimBus9[6];
assign
s_logisimBus21[8]
=
s_logisimBus9[7];
assign
s_logisimBus21[9]
=
s_logisimBus9[8];
assign
s_logisimBus34[0]
=
s_logisimBus6[0];
assign
s_logisimBus34[10]
=
s_logisimBus6[10];
assign
s_logisimBus34[11]
=
s_logisimBus6[11];
assign
s_logisimBus34[12]
=
s_logisimBus6[12];
assign
s_logisimBus34[13]
=
s_logisimBus6[13];
assign
s_logisimBus34[14]
=
s_logisimBus6[14];
assign
s_logisimBus34[15]
=
s_logisimBus6[15];
assign
s_logisimBus34[16]
=
s_logisimBus6[16];
assign
s_logisimBus34[17]
=
s_logisimBus6[17];
assign
s_logisimBus34[18]
=
s_logisimBus6[18];
assign
s_logisimBus34[19]
=
s_logisimBus6[19];
assign
s_logisimBus34[1]
=
s_logisimBus6[1];
assign
s_logisimBus34[20]
=
s_logisimBus6[20];
assign
s_logisimBus34[21]
=
s_logisimBus6[21];
assign
s_logisimBus34[22]
=
s_logisimBus6[22];
assign
s_logisimBus34[23]
=
s_logisimBus6[23];
assign
s_logisimBus34[24]
=
s_logisimBus6[24];
assign
s_logisimBus34[25]
=
s_logisimBus6[25];
assign
s_logisimBus34[26]
=
s_logisimBus6[26];
assign
s_logisimBus34[27]
=
s_logisimBus6[27];
assign
s_logisimBus34[28]
=
s_logisimBus6[28];
assign
s_logisimBus34[29]
=
s_logisimBus6[29];
assign
s_logisimBus34[2]
=
s_logisimBus6[2];
assign
s_logisimBus34[30]
=
s_logisimBus6[30];
assign
s_logisimBus34[3]
=
s_logisimBus6[3];
assign
s_logisimBus34[4]
=
s_logisimBus6[4];
assign
s_logisimBus34[5]
=
s_logisimBus6[5];
assign
s_logisimBus34[6]
=
s_logisimBus6[6];
assign
s_logisimBus34[7]
=
s_logisimBus6[7];
assign
s_logisimBus34[8]
=
s_logisimBus6[8];
assign
s_logisimBus34[9]
=
s_logisimBus6[9];
assign
s_logisimBus4[0]
=
s_logisimNet23;
assign
s_logisimBus4[10]
=
s_logisimBus34[9];
assign
s_logisimBus4[11]
=
s_logisimBus34[10];
assign
s_logisimBus4[12]
=
s_logisimBus34[11];
assign
s_logisimBus4[13]
=
s_logisimBus34[12];
assign
s_logisimBus4[14]
=
s_logisimBus34[13];
assign
s_logisimBus4[15]
=
s_logisimBus34[14];
assign
s_logisimBus4[16]
=
s_logisimBus34[15];
assign
s_logisimBus4[17]
=
s_logisimBus34[16];
assign
s_logisimBus4[18]
=
s_logisimBus34[17];
assign
s_logisimBus4[19]
=
s_logisimBus34[18];
assign
s_logisimBus4[1]
=
s_logisimBus34[0];
assign
s_logisimBus4[20]
=
s_logisimBus34[19];
assign
s_logisimBus4[21]
=
s_logisimBus34[20];
assign
s_logisimBus4[22]
=
s_logisimBus34[21];
assign
s_logisimBus4[23]
=
s_logisimBus34[22];
assign
s_logisimBus4[24]
=
s_logisimBus34[23];
assign
s_logisimBus4[25]
=
s_logisimBus34[24];
assign
s_logisimBus4[26]
=
s_logisimBus34[25];
assign
s_logisimBus4[27]
=
s_logisimBus34[26];
assign
s_logisimBus4[28]
=
s_logisimBus34[27];
assign
s_logisimBus4[29]
=
s_logisimBus34[28];
assign
s_logisimBus4[2]
=
s_logisimBus34[1];
assign
s_logisimBus4[30]
=
s_logisimBus34[29];
assign
s_logisimBus4[31]
=
s_logisimBus34[30];
assign
s_logisimBus4[3]
=
s_logisimBus34[2];
assign
s_logisimBus4[4]
=
s_logisimBus34[3];
assign
s_logisimBus4[5]
=
s_logisimBus34[4];
assign
s_logisimBus4[6]
=
s_logisimBus34[5];
assign
s_logisimBus4[7]
=
s_logisimBus34[6];
assign
s_logisimBus4[8]
=
s_logisimBus34[7];
assign
s_logisimBus4[9]
=
s_logisimBus34[8];
assign
s_logisimBus9[0]
=
s_logisimBus32[0];
assign
s_logisimBus9[10]
=
s_logisimBus32[10];
assign
s_logisimBus9[11]
=
s_logisimBus32[11];
assign
s_logisimBus9[12]
=
s_logisimBus32[12];
assign
s_logisimBus9[13]
=
s_logisimBus32[13];
assign
s_logisimBus9[14]
=
s_logisimBus32[14];
assign
s_logisimBus9[15]
=
s_logisimBus32[15];
assign
s_logisimBus9[16]
=
s_logisimBus32[16];
assign
s_logisimBus9[17]
=
s_logisimBus32[17];
assign
s_logisimBus9[18]
=
s_logisimBus32[18];
assign
s_logisimBus9[19]
=
s_logisimBus32[19];
assign
s_logisimBus9[1]
=
s_logisimBus32[1];
assign
s_logisimBus9[20]
=
s_logisimBus32[20];
assign
s_logisimBus9[21]
=
s_logisimBus32[21];
assign
s_logisimBus9[22]
=
s_logisimBus32[22];
assign
s_logisimBus9[23]
=
s_logisimBus32[23];
assign
s_logisimBus9[24]
=
s_logisimBus32[24];
assign
s_logisimBus9[25]
=
s_logisimBus32[25];
assign
s_logisimBus9[26]
=
s_logisimBus32[26];
assign
s_logisimBus9[27]
=
s_logisimBus32[27];
assign
s_logisimBus9[28]
=
s_logisimBus32[28];
assign
s_logisimBus9[29]
=
s_logisimBus32[29];
assign
s_logisimBus9[2]
=
s_logisimBus32[2];
assign
s_logisimBus9[30]
=
s_logisimBus32[30];
assign
s_logisimBus9[3]
=
s_logisimBus32[3];
assign
s_logisimBus9[4]
=
s_logisimBus32[4];
assign
s_logisimBus9[5]
=
s_logisimBus32[5];
assign
s_logisimBus9[6]
=
s_logisimBus32[6];
assign
s_logisimBus9[7]
=
s_logisimBus32[7];
assign
s_logisimBus9[8]
=
s_logisimBus32[8];
assign
s_logisimBus9[9]
=
s_logisimBus32[9];
assign
s_logisimNet23
=
s_logisimBus32[31];
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus1[31:0]
=
divisor;
assign
s_logisimBus27[31:0]
=
dividend;
assign
s_logisimNet8
=
clk;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
done
=
s_logisimNet11;
assign
quotient
=
s_logisimBus19[31:0];
assign
remainder
=
s_logisimBus20[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimNet38
=
1'b1;
assign
s_logisimNet39
=
1'b1;
assign
s_logisimBus28[63:0]
=
64'h0000000000000020;
assign
s_logisimNet37
=
1'b1;
assign
s_logisimNet30
=
1'b0;
assign
s_logisimNet22
=
1'b1;
assign
s_logisimNet33
=
1'b1;
assign
s_logisimNet14
=
1'b0;
assign
s_logisimBus5[63:0]
=
64'h0000000000000000;
assign
s_logisimBus29[63:0]
=
64'h0000000000000001;
assign
s_logisimNet7
=
1'b0;
assign
s_logisimNet24
=
1'b0;
assign
s_logisimNet17
=
~s_logisimNet31;
assign
s_logisimNet12
=
~s_logisimNet15;
assign
s_logisimBus21[0]
=
~s_logisimNet16;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE
#(.BubblesMask(2'b00))
GATES_1
(.input1(s_logisimNet17),
.input2(s_logisimNet12),
.result(s_logisimNet2));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus25[63:0]),
.muxIn_1(s_logisimBus28[63:0]),
.muxOut(s_logisimBus35[63:0]),
.sel(s_logisimNet2));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus21[31:0]),
.muxIn_1(s_logisimBus27[31:0]),
.muxOut(s_logisimBus10[31:0]),
.sel(s_logisimNet2));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus3[31:0]),
.muxIn_1(s_logisimBus36[31:0]),
.muxOut(s_logisimBus6[31:0]),
.sel(s_logisimBus21[0]));
Comparator
#(.nrOfBits(32),
.twosComplement(0))
ARITH_5
(.aEqualsB(s_logisimNet31),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus27[31:0]),
.dataB(s_logisimBus13[31:0]));
Comparator
#(.nrOfBits(32),
.twosComplement(0))
ARITH_6
(.aEqualsB(s_logisimNet15),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus1[31:0]),
.dataB(s_logisimBus18[31:0]));
Subtractor
#(.extendedBits(33),
.nrOfBits(32))
ARITH_7
(.borrowIn(s_logisimNet7),
.borrowOut(),
.dataA(s_logisimBus3[31:0]),
.dataB(s_logisimBus1[31:0]),
.result(s_logisimBus36[31:0]));
Comparator
#(.nrOfBits(32),
.twosComplement(0))
ARITH_8
(.aEqualsB(),
.aGreaterThanB(),
.aLessThanB(s_logisimNet16),
.dataA(s_logisimBus3[31:0]),
.dataB(s_logisimBus1[31:0]));
Subtractor
#(.extendedBits(65),
.nrOfBits(64))
ARITH_9
(.borrowIn(s_logisimNet24),
.borrowOut(),
.dataA(s_logisimBus0[63:0]),
.dataB(s_logisimBus29[63:0]),
.result(s_logisimBus25[63:0]));
Comparator
#(.nrOfBits(64),
.twosComplement(0))
ARITH_10
(.aEqualsB(s_logisimNet11),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus0[63:0]),
.dataB(s_logisimBus5[63:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_11
(.clock(s_logisimNet8),
.clockEnable(s_logisimNet38),
.d(s_logisimBus27[31:0]),
.q(s_logisimBus13[31:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_12
(.clock(s_logisimNet8),
.clockEnable(s_logisimNet39),
.d(s_logisimBus1[31:0]),
.q(s_logisimBus18[31:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(64))
counter
(.clock(s_logisimNet8),
.clockEnable(s_logisimNet37),
.d(s_logisimBus35[63:0]),
.q(s_logisimBus0[63:0]),
.reset(s_logisimNet30),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
q_reg
(.clock(s_logisimNet8),
.clockEnable(s_logisimNet22),
.d(s_logisimBus10[31:0]),
.q(s_logisimBus32[31:0]),
.reset(s_logisimNet14),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
a_reg
(.clock(s_logisimNet8),
.clockEnable(s_logisimNet33),
.d(s_logisimBus4[31:0]),
.q(s_logisimBus3[31:0]),
.reset(s_logisimNet2),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_16
(.clock(s_logisimNet8),
.clockEnable(s_logisimNet11),
.d(s_logisimBus21[31:0]),
.q(s_logisimBus19[31:0]),
.reset(s_logisimNet2),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_17
(.clock(s_logisimNet8),
.clockEnable(s_logisimNet11),
.d(s_logisimBus6[31:0]),
.q(s_logisimBus20[31:0]),
.reset(s_logisimNet2),
.tick(1'b1));
endmodule