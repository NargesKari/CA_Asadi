/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
SRA11
**
**
**
*****************************************************************************/
module
SRA11(
a,
b,
output1
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[31:0]
b;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[63:0]
output1;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[63:0]
s_logisimBus10;
wire
[31:0]
s_logisimBus12;
wire
[63:0]
s_logisimBus13;
wire
[63:0]
s_logisimBus14;
wire
[5:0]
s_logisimBus16;
wire
[63:0]
s_logisimBus17;
wire
[31:0]
s_logisimBus20;
wire
[31:0]
s_logisimBus22;
wire
[5:0]
s_logisimBus24;
wire
[31:0]
s_logisimBus25;
wire
[63:0]
s_logisimBus26;
wire
[31:0]
s_logisimBus27;
wire
[31:0]
s_logisimBus3;
wire
[31:0]
s_logisimBus4;
wire
[7:0]
s_logisimBus5;
wire
[63:0]
s_logisimBus6;
wire
[63:0]
s_logisimBus7;
wire
[31:0]
s_logisimBus8;
wire
[31:0]
s_logisimBus9;
wire
s_logisimNet15;
wire
s_logisimNet18;
wire
s_logisimNet23;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
wiring
is
defined
**
*******************************************************************************/
assign
s_logisimBus10[0]
=
s_logisimBus8[0];
assign
s_logisimBus10[10]
=
s_logisimBus8[10];
assign
s_logisimBus10[11]
=
s_logisimBus8[11];
assign
s_logisimBus10[12]
=
s_logisimBus8[12];
assign
s_logisimBus10[13]
=
s_logisimBus8[13];
assign
s_logisimBus10[14]
=
s_logisimBus8[14];
assign
s_logisimBus10[15]
=
s_logisimBus8[15];
assign
s_logisimBus10[16]
=
s_logisimBus8[16];
assign
s_logisimBus10[17]
=
s_logisimBus8[17];
assign
s_logisimBus10[18]
=
s_logisimBus8[18];
assign
s_logisimBus10[19]
=
s_logisimBus8[19];
assign
s_logisimBus10[1]
=
s_logisimBus8[1];
assign
s_logisimBus10[20]
=
s_logisimBus8[20];
assign
s_logisimBus10[21]
=
s_logisimBus8[21];
assign
s_logisimBus10[22]
=
s_logisimBus8[22];
assign
s_logisimBus10[23]
=
s_logisimBus8[23];
assign
s_logisimBus10[24]
=
s_logisimBus8[24];
assign
s_logisimBus10[25]
=
s_logisimBus8[25];
assign
s_logisimBus10[26]
=
s_logisimBus8[26];
assign
s_logisimBus10[27]
=
s_logisimBus8[27];
assign
s_logisimBus10[28]
=
s_logisimBus8[28];
assign
s_logisimBus10[29]
=
s_logisimBus8[29];
assign
s_logisimBus10[2]
=
s_logisimBus8[2];
assign
s_logisimBus10[30]
=
s_logisimBus8[30];
assign
s_logisimBus10[31]
=
s_logisimBus8[31];
assign
s_logisimBus10[3]
=
s_logisimBus8[3];
assign
s_logisimBus10[4]
=
s_logisimBus8[4];
assign
s_logisimBus10[5]
=
s_logisimBus8[5];
assign
s_logisimBus10[6]
=
s_logisimBus8[6];
assign
s_logisimBus10[7]
=
s_logisimBus8[7];
assign
s_logisimBus10[8]
=
s_logisimBus8[8];
assign
s_logisimBus10[9]
=
s_logisimBus8[9];
assign
s_logisimBus4[16]
=
s_logisimBus5[0];
assign
s_logisimBus4[17]
=
s_logisimBus5[1];
assign
s_logisimBus4[18]
=
s_logisimBus5[2];
assign
s_logisimBus4[19]
=
s_logisimBus5[3];
assign
s_logisimBus4[20]
=
s_logisimBus5[4];
assign
s_logisimBus4[21]
=
s_logisimBus5[5];
assign
s_logisimBus4[22]
=
s_logisimBus5[6];
assign
s_logisimBus4[23]
=
s_logisimBus5[7];
assign
s_logisimBus4[24]
=
s_logisimBus5[0];
assign
s_logisimBus4[25]
=
s_logisimBus5[1];
assign
s_logisimBus4[26]
=
s_logisimBus5[2];
assign
s_logisimBus4[27]
=
s_logisimBus5[3];
assign
s_logisimBus4[28]
=
s_logisimBus5[4];
assign
s_logisimBus4[29]
=
s_logisimBus5[5];
assign
s_logisimBus4[30]
=
s_logisimBus5[6];
assign
s_logisimBus4[31]
=
s_logisimBus5[7];
assign
s_logisimBus8[0]
=
s_logisimBus13[0];
assign
s_logisimBus8[10]
=
s_logisimBus13[10];
assign
s_logisimBus8[11]
=
s_logisimBus13[11];
assign
s_logisimBus8[12]
=
s_logisimBus13[12];
assign
s_logisimBus8[13]
=
s_logisimBus13[13];
assign
s_logisimBus8[14]
=
s_logisimBus13[14];
assign
s_logisimBus8[15]
=
s_logisimBus13[15];
assign
s_logisimBus8[16]
=
s_logisimBus13[16];
assign
s_logisimBus8[17]
=
s_logisimBus13[17];
assign
s_logisimBus8[18]
=
s_logisimBus13[18];
assign
s_logisimBus8[19]
=
s_logisimBus13[19];
assign
s_logisimBus8[1]
=
s_logisimBus13[1];
assign
s_logisimBus8[20]
=
s_logisimBus13[20];
assign
s_logisimBus8[21]
=
s_logisimBus13[21];
assign
s_logisimBus8[22]
=
s_logisimBus13[22];
assign
s_logisimBus8[23]
=
s_logisimBus13[23];
assign
s_logisimBus8[24]
=
s_logisimBus13[24];
assign
s_logisimBus8[25]
=
s_logisimBus13[25];
assign
s_logisimBus8[26]
=
s_logisimBus13[26];
assign
s_logisimBus8[27]
=
s_logisimBus13[27];
assign
s_logisimBus8[28]
=
s_logisimBus13[28];
assign
s_logisimBus8[29]
=
s_logisimBus13[29];
assign
s_logisimBus8[2]
=
s_logisimBus13[2];
assign
s_logisimBus8[30]
=
s_logisimBus13[30];
assign
s_logisimBus8[31]
=
s_logisimBus13[31];
assign
s_logisimBus8[3]
=
s_logisimBus13[3];
assign
s_logisimBus8[4]
=
s_logisimBus13[4];
assign
s_logisimBus8[5]
=
s_logisimBus13[5];
assign
s_logisimBus8[6]
=
s_logisimBus13[6];
assign
s_logisimBus8[7]
=
s_logisimBus13[7];
assign
s_logisimBus8[8]
=
s_logisimBus13[8];
assign
s_logisimBus8[9]
=
s_logisimBus13[9];
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus12[31:0]
=
a;
assign
s_logisimBus27[31:0]
=
b;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
output1
=
s_logisimBus10[63:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus5[7:0]
=
8'h00;
assign
s_logisimBus4[0]
=
s_logisimBus27[0];
assign
s_logisimBus4[1]
=
s_logisimBus27[1];
assign
s_logisimBus4[2]
=
s_logisimBus27[2];
assign
s_logisimBus4[3]
=
s_logisimBus27[3];
assign
s_logisimBus4[4]
=
s_logisimBus27[4];
assign
s_logisimBus7[0]
=
s_logisimBus12[0];
assign
s_logisimBus7[1]
=
s_logisimBus12[1];
assign
s_logisimBus7[2]
=
s_logisimBus12[2];
assign
s_logisimBus7[3]
=
s_logisimBus12[3];
assign
s_logisimBus7[4]
=
s_logisimBus12[4];
assign
s_logisimBus7[5]
=
s_logisimBus12[5];
assign
s_logisimBus7[6]
=
s_logisimBus12[6];
assign
s_logisimBus7[7]
=
s_logisimBus12[7];
assign
s_logisimBus7[8]
=
s_logisimBus12[8];
assign
s_logisimBus7[9]
=
s_logisimBus12[9];
assign
s_logisimBus7[10]
=
s_logisimBus12[10];
assign
s_logisimBus7[11]
=
s_logisimBus12[11];
assign
s_logisimBus7[12]
=
s_logisimBus12[12];
assign
s_logisimBus7[13]
=
s_logisimBus12[13];
assign
s_logisimBus7[14]
=
s_logisimBus12[14];
assign
s_logisimBus7[15]
=
s_logisimBus12[15];
assign
s_logisimBus7[16]
=
s_logisimBus12[16];
assign
s_logisimBus7[17]
=
s_logisimBus12[17];
assign
s_logisimBus7[18]
=
s_logisimBus12[18];
assign
s_logisimBus7[19]
=
s_logisimBus12[19];
assign
s_logisimBus7[20]
=
s_logisimBus12[20];
assign
s_logisimBus7[21]
=
s_logisimBus12[21];
assign
s_logisimBus7[22]
=
s_logisimBus12[22];
assign
s_logisimBus7[23]
=
s_logisimBus12[23];
assign
s_logisimBus7[24]
=
s_logisimBus12[24];
assign
s_logisimBus7[25]
=
s_logisimBus12[25];
assign
s_logisimBus7[26]
=
s_logisimBus12[26];
assign
s_logisimBus7[27]
=
s_logisimBus12[27];
assign
s_logisimBus7[28]
=
s_logisimBus12[28];
assign
s_logisimBus7[29]
=
s_logisimBus12[29];
assign
s_logisimBus7[30]
=
s_logisimBus12[30];
assign
s_logisimBus7[31]
=
s_logisimBus12[31];
assign
s_logisimBus7[32]
=
s_logisimBus12[31];
assign
s_logisimBus7[33]
=
s_logisimBus12[31];
assign
s_logisimBus7[34]
=
s_logisimBus12[31];
assign
s_logisimBus7[35]
=
s_logisimBus12[31];
assign
s_logisimBus7[36]
=
s_logisimBus12[31];
assign
s_logisimBus7[37]
=
s_logisimBus12[31];
assign
s_logisimBus7[38]
=
s_logisimBus12[31];
assign
s_logisimBus7[39]
=
s_logisimBus12[31];
assign
s_logisimBus7[40]
=
s_logisimBus12[31];
assign
s_logisimBus7[41]
=
s_logisimBus12[31];
assign
s_logisimBus7[42]
=
s_logisimBus12[31];
assign
s_logisimBus7[43]
=
s_logisimBus12[31];
assign
s_logisimBus7[44]
=
s_logisimBus12[31];
assign
s_logisimBus7[45]
=
s_logisimBus12[31];
assign
s_logisimBus7[46]
=
s_logisimBus12[31];
assign
s_logisimBus7[47]
=
s_logisimBus12[31];
assign
s_logisimBus7[48]
=
s_logisimBus12[31];
assign
s_logisimBus7[49]
=
s_logisimBus12[31];
assign
s_logisimBus7[50]
=
s_logisimBus12[31];
assign
s_logisimBus7[51]
=
s_logisimBus12[31];
assign
s_logisimBus7[52]
=
s_logisimBus12[31];
assign
s_logisimBus7[53]
=
s_logisimBus12[31];
assign
s_logisimBus7[54]
=
s_logisimBus12[31];
assign
s_logisimBus7[55]
=
s_logisimBus12[31];
assign
s_logisimBus7[56]
=
s_logisimBus12[31];
assign
s_logisimBus7[57]
=
s_logisimBus12[31];
assign
s_logisimBus7[58]
=
s_logisimBus12[31];
assign
s_logisimBus7[59]
=
s_logisimBus12[31];
assign
s_logisimBus7[60]
=
s_logisimBus12[31];
assign
s_logisimBus7[61]
=
s_logisimBus12[31];
assign
s_logisimBus7[62]
=
s_logisimBus12[31];
assign
s_logisimBus7[63]
=
s_logisimBus12[31];
assign
s_logisimBus16[5:0]
=
{2'b00,
4'h1};
assign
s_logisimBus22[31:0]
=
32'h00000001;
assign
s_logisimBus4[15:5]
=
{3'b000,
8'h00};
assign
s_logisimBus24[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus20[31:0]
=
32'h00000000;
assign
s_logisimBus0[31:0]
=
32'hFFFFFFFF;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_1
(.enable(1'b1),
.muxIn_0(s_logisimBus14[63:0]),
.muxIn_1(s_logisimBus26[63:0]),
.muxOut(s_logisimBus17[63:0]),
.sel(s_logisimBus4[0]));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus20[31:0]),
.muxIn_1(s_logisimBus0[31:0]),
.muxOut(s_logisimBus10[63:32]),
.sel(s_logisimBus13[31]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus17[63:0]),
.muxIn_1(s_logisimBus7[63:0]),
.muxOut(s_logisimBus13[63:0]),
.sel(s_logisimNet15));
Shifter_64_bit
#(.shifterMode(2))
ARITH_4
(.dataA(s_logisimBus7[63:0]),
.result(s_logisimBus6[63:0]),
.shiftAmount(s_logisimBus16[5:0]));
Subtractor
#(.extendedBits(33),
.nrOfBits(32))
ARITH_5
(.borrowIn(1'b0),
.borrowOut(),
.dataA(s_logisimBus4[31:0]),
.dataB(s_logisimBus22[31:0]),
.result(s_logisimBus25[31:0]));
Shifter_64_bit
#(.shifterMode(2))
ARITH_6
(.dataA(s_logisimBus7[63:0]),
.result(s_logisimBus26[63:0]),
.shiftAmount(s_logisimBus4[5:0]));
Shifter_64_bit
#(.shifterMode(2))
ARITH_7
(.dataA(s_logisimBus6[63:0]),
.result(s_logisimBus14[63:0]),
.shiftAmount(s_logisimBus25[5:0]));
Comparator
#(.nrOfBits(32),
.twosComplement(1))
ARITH_8
(.aEqualsB(),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[31:0]),
.dataB(s_logisimBus3[31:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_9
(.aEqualsB(s_logisimNet15),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus4[5:0]),
.dataB(s_logisimBus24[5:0]));
endmodule