/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
ALU_CLO
**
**
**
*****************************************************************************/
module
ALU_CLO(
A,
OUTTTT
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
A;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[63:0]
OUTTTT;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[3:0]
s_logisimBus100;
wire
[3:0]
s_logisimBus102;
wire
[2:0]
s_logisimBus103;
wire
[63:0]
s_logisimBus105;
wire
[1:0]
s_logisimBus114;
wire
[1:0]
s_logisimBus115;
wire
[1:0]
s_logisimBus116;
wire
[1:0]
s_logisimBus117;
wire
[63:0]
s_logisimBus12;
wire
[1:0]
s_logisimBus2;
wire
[2:0]
s_logisimBus35;
wire
[2:0]
s_logisimBus47;
wire
[2:0]
s_logisimBus64;
wire
[63:0]
s_logisimBus78;
wire
[1:0]
s_logisimBus81;
wire
[1:0]
s_logisimBus92;
wire
[1:0]
s_logisimBus95;
wire
[31:0]
s_logisimBus99;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet101;
wire
s_logisimNet104;
wire
s_logisimNet106;
wire
s_logisimNet107;
wire
s_logisimNet109;
wire
s_logisimNet11;
wire
s_logisimNet112;
wire
s_logisimNet113;
wire
s_logisimNet13;
wire
s_logisimNet14;
wire
s_logisimNet16;
wire
s_logisimNet17;
wire
s_logisimNet18;
wire
s_logisimNet19;
wire
s_logisimNet20;
wire
s_logisimNet21;
wire
s_logisimNet22;
wire
s_logisimNet25;
wire
s_logisimNet26;
wire
s_logisimNet27;
wire
s_logisimNet28;
wire
s_logisimNet29;
wire
s_logisimNet3;
wire
s_logisimNet30;
wire
s_logisimNet32;
wire
s_logisimNet33;
wire
s_logisimNet34;
wire
s_logisimNet36;
wire
s_logisimNet37;
wire
s_logisimNet38;
wire
s_logisimNet39;
wire
s_logisimNet4;
wire
s_logisimNet40;
wire
s_logisimNet41;
wire
s_logisimNet42;
wire
s_logisimNet43;
wire
s_logisimNet44;
wire
s_logisimNet45;
wire
s_logisimNet46;
wire
s_logisimNet48;
wire
s_logisimNet49;
wire
s_logisimNet5;
wire
s_logisimNet50;
wire
s_logisimNet51;
wire
s_logisimNet52;
wire
s_logisimNet54;
wire
s_logisimNet55;
wire
s_logisimNet56;
wire
s_logisimNet57;
wire
s_logisimNet58;
wire
s_logisimNet59;
wire
s_logisimNet6;
wire
s_logisimNet60;
wire
s_logisimNet61;
wire
s_logisimNet62;
wire
s_logisimNet63;
wire
s_logisimNet65;
wire
s_logisimNet66;
wire
s_logisimNet67;
wire
s_logisimNet68;
wire
s_logisimNet69;
wire
s_logisimNet7;
wire
s_logisimNet70;
wire
s_logisimNet71;
wire
s_logisimNet73;
wire
s_logisimNet74;
wire
s_logisimNet75;
wire
s_logisimNet76;
wire
s_logisimNet77;
wire
s_logisimNet79;
wire
s_logisimNet8;
wire
s_logisimNet82;
wire
s_logisimNet83;
wire
s_logisimNet84;
wire
s_logisimNet85;
wire
s_logisimNet86;
wire
s_logisimNet87;
wire
s_logisimNet88;
wire
s_logisimNet89;
wire
s_logisimNet9;
wire
s_logisimNet90;
wire
s_logisimNet91;
wire
s_logisimNet93;
wire
s_logisimNet94;
wire
s_logisimNet96;
wire
s_logisimNet97;
wire
s_logisimNet98;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus99[31:0]
=
A;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
OUTTTT
=
s_logisimBus105[63:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus12[52:37]
=
16'h0000;
assign
s_logisimBus12[62:61]
=
2'b00;
assign
s_logisimBus78[63:0]
=
64'h0000000000000000;
assign
s_logisimBus12[60:53]
=
8'h00;
assign
s_logisimBus12[36:5]
=
32'h00000000;
assign
s_logisimBus12[63]
=
1'b0;
assign
s_logisimNet75
=
1'b1;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE
#(.BubblesMask(2'b00))
GATES_1
(.input1(s_logisimBus99[16]),
.input2(s_logisimNet89),
.result(s_logisimNet48));
AND_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimBus99[15]),
.input2(s_logisimNet48),
.result(s_logisimNet11));
AND_GATE
#(.BubblesMask(2'b00))
GATES_3
(.input1(s_logisimBus99[14]),
.input2(s_logisimNet11),
.result(s_logisimNet25));
AND_GATE
#(.BubblesMask(2'b00))
GATES_4
(.input1(s_logisimBus99[13]),
.input2(s_logisimNet25),
.result(s_logisimNet76));
AND_GATE
#(.BubblesMask(2'b00))
GATES_5
(.input1(s_logisimBus99[12]),
.input2(s_logisimNet76),
.result(s_logisimNet7));
AND_GATE
#(.BubblesMask(2'b00))
GATES_6
(.input1(s_logisimBus99[11]),
.input2(s_logisimNet7),
.result(s_logisimNet9));
AND_GATE
#(.BubblesMask(2'b00))
GATES_7
(.input1(s_logisimBus99[10]),
.input2(s_logisimNet9),
.result(s_logisimNet56));
AND_GATE
#(.BubblesMask(2'b00))
GATES_8
(.input1(s_logisimBus99[9]),
.input2(s_logisimNet56),
.result(s_logisimNet8));
AND_GATE
#(.BubblesMask(2'b00))
GATES_9
(.input1(s_logisimBus99[8]),
.input2(s_logisimNet8),
.result(s_logisimNet39));
AND_GATE
#(.BubblesMask(2'b00))
GATES_10
(.input1(s_logisimBus99[7]),
.input2(s_logisimNet39),
.result(s_logisimNet5));
AND_GATE
#(.BubblesMask(2'b00))
GATES_11
(.input1(s_logisimBus99[6]),
.input2(s_logisimNet5),
.result(s_logisimNet50));
AND_GATE
#(.BubblesMask(2'b00))
GATES_12
(.input1(s_logisimBus99[5]),
.input2(s_logisimNet50),
.result(s_logisimNet66));
AND_GATE
#(.BubblesMask(2'b00))
GATES_13
(.input1(s_logisimBus99[4]),
.input2(s_logisimNet66),
.result(s_logisimNet30));
AND_GATE
#(.BubblesMask(2'b00))
GATES_14
(.input1(s_logisimBus99[3]),
.input2(s_logisimNet30),
.result(s_logisimNet6));
AND_GATE
#(.BubblesMask(2'b00))
GATES_15
(.input1(s_logisimBus99[2]),
.input2(s_logisimNet6),
.result(s_logisimNet58));
AND_GATE
#(.BubblesMask(2'b00))
GATES_16
(.input1(s_logisimBus99[1]),
.input2(s_logisimNet58),
.result(s_logisimNet17));
AND_GATE
#(.BubblesMask(2'b00))
GATES_17
(.input1(s_logisimBus99[0]),
.input2(s_logisimNet17),
.result(s_logisimNet13));
AND_GATE
#(.BubblesMask(2'b00))
GATES_18
(.input1(s_logisimBus99[31]),
.input2(s_logisimNet75),
.result(s_logisimNet18));
AND_GATE
#(.BubblesMask(2'b00))
GATES_19
(.input1(s_logisimBus99[30]),
.input2(s_logisimNet18),
.result(s_logisimNet28));
AND_GATE
#(.BubblesMask(2'b00))
GATES_20
(.input1(s_logisimBus99[29]),
.input2(s_logisimNet28),
.result(s_logisimNet69));
AND_GATE
#(.BubblesMask(2'b00))
GATES_21
(.input1(s_logisimBus99[28]),
.input2(s_logisimNet69),
.result(s_logisimNet44));
AND_GATE
#(.BubblesMask(2'b00))
GATES_22
(.input1(s_logisimBus99[27]),
.input2(s_logisimNet44),
.result(s_logisimNet16));
AND_GATE
#(.BubblesMask(2'b00))
GATES_23
(.input1(s_logisimBus99[26]),
.input2(s_logisimNet16),
.result(s_logisimNet34));
AND_GATE
#(.BubblesMask(2'b00))
GATES_24
(.input1(s_logisimBus99[25]),
.input2(s_logisimNet34),
.result(s_logisimNet88));
AND_GATE
#(.BubblesMask(2'b00))
GATES_25
(.input1(s_logisimBus99[24]),
.input2(s_logisimNet88),
.result(s_logisimNet51));
AND_GATE
#(.BubblesMask(2'b00))
GATES_26
(.input1(s_logisimBus99[23]),
.input2(s_logisimNet51),
.result(s_logisimNet22));
AND_GATE
#(.BubblesMask(2'b00))
GATES_27
(.input1(s_logisimBus99[22]),
.input2(s_logisimNet22),
.result(s_logisimNet36));
AND_GATE
#(.BubblesMask(2'b00))
GATES_28
(.input1(s_logisimBus99[21]),
.input2(s_logisimNet36),
.result(s_logisimNet73));
AND_GATE
#(.BubblesMask(2'b00))
GATES_29
(.input1(s_logisimBus99[20]),
.input2(s_logisimNet73),
.result(s_logisimNet20));
AND_GATE
#(.BubblesMask(2'b00))
GATES_30
(.input1(s_logisimBus99[19]),
.input2(s_logisimNet20),
.result(s_logisimNet21));
AND_GATE
#(.BubblesMask(2'b00))
GATES_31
(.input1(s_logisimBus99[18]),
.input2(s_logisimNet21),
.result(s_logisimNet60));
AND_GATE
#(.BubblesMask(2'b00))
GATES_32
(.input1(s_logisimBus99[17]),
.input2(s_logisimNet60),
.result(s_logisimNet89));
FullAdder
#(.extendedBits(2))
ARITH_33
(.carryIn(s_logisimNet25),
.carryOut(s_logisimBus95[1]),
.dataA(s_logisimNet11),
.dataB(s_logisimNet48),
.result(s_logisimBus95[0]));
FullAdder
#(.extendedBits(2))
ARITH_34
(.carryIn(s_logisimNet9),
.carryOut(s_logisimBus114[1]),
.dataA(s_logisimNet7),
.dataB(s_logisimNet76),
.result(s_logisimBus114[0]));
Adder
#(.extendedBits(3),
.nrOfBits(2))
ARITH_35
(.carryIn(s_logisimNet56),
.carryOut(s_logisimBus35[2]),
.dataA(s_logisimBus114[1:0]),
.dataB(s_logisimBus95[1:0]),
.result(s_logisimBus35[1:0]));
FullAdder
#(.extendedBits(2))
ARITH_36
(.carryIn(s_logisimNet5),
.carryOut(s_logisimBus81[1]),
.dataA(s_logisimNet39),
.dataB(s_logisimNet8),
.result(s_logisimBus81[0]));
FullAdder
#(.extendedBits(2))
ARITH_37
(.carryIn(s_logisimNet30),
.carryOut(s_logisimBus115[1]),
.dataA(s_logisimNet66),
.dataB(s_logisimNet50),
.result(s_logisimBus115[0]));
Adder
#(.extendedBits(3),
.nrOfBits(2))
ARITH_38
(.carryIn(s_logisimNet6),
.carryOut(s_logisimBus103[2]),
.dataA(s_logisimBus115[1:0]),
.dataB(s_logisimBus81[1:0]),
.result(s_logisimBus103[1:0]));
Adder
#(.extendedBits(4),
.nrOfBits(3))
ARITH_39
(.carryIn(s_logisimNet58),
.carryOut(s_logisimBus102[3]),
.dataA(s_logisimBus103[2:0]),
.dataB(s_logisimBus35[2:0]),
.result(s_logisimBus102[2:0]));
Adder
#(.extendedBits(5),
.nrOfBits(4))
ARITH_40
(.carryIn(s_logisimNet17),
.carryOut(s_logisimBus12[4]),
.dataA(s_logisimBus102[3:0]),
.dataB(s_logisimBus100[3:0]),
.result(s_logisimBus12[3:0]));
Adder
#(.extendedBits(65),
.nrOfBits(64))
ARITH_41
(.carryIn(s_logisimNet13),
.carryOut(),
.dataA(s_logisimBus78[63:0]),
.dataB(s_logisimBus12[63:0]),
.result(s_logisimBus105[63:0]));
FullAdder
#(.extendedBits(2))
ARITH_42
(.carryIn(s_logisimNet69),
.carryOut(s_logisimBus2[1]),
.dataA(s_logisimNet28),
.dataB(s_logisimNet18),
.result(s_logisimBus2[0]));
FullAdder
#(.extendedBits(2))
ARITH_43
(.carryIn(s_logisimNet34),
.carryOut(s_logisimBus116[1]),
.dataA(s_logisimNet16),
.dataB(s_logisimNet44),
.result(s_logisimBus116[0]));
Adder
#(.extendedBits(3),
.nrOfBits(2))
ARITH_44
(.carryIn(s_logisimNet88),
.carryOut(s_logisimBus64[2]),
.dataA(s_logisimBus116[1:0]),
.dataB(s_logisimBus2[1:0]),
.result(s_logisimBus64[1:0]));
FullAdder
#(.extendedBits(2))
ARITH_45
(.carryIn(s_logisimNet36),
.carryOut(s_logisimBus92[1]),
.dataA(s_logisimNet22),
.dataB(s_logisimNet51),
.result(s_logisimBus92[0]));
FullAdder
#(.extendedBits(2))
ARITH_46
(.carryIn(s_logisimNet21),
.carryOut(s_logisimBus117[1]),
.dataA(s_logisimNet20),
.dataB(s_logisimNet73),
.result(s_logisimBus117[0]));
Adder
#(.extendedBits(3),
.nrOfBits(2))
ARITH_47
(.carryIn(s_logisimNet60),
.carryOut(s_logisimBus47[2]),
.dataA(s_logisimBus117[1:0]),
.dataB(s_logisimBus92[1:0]),
.result(s_logisimBus47[1:0]));
Adder
#(.extendedBits(4),
.nrOfBits(3))
ARITH_48
(.carryIn(s_logisimNet89),
.carryOut(s_logisimBus100[3]),
.dataA(s_logisimBus47[2:0]),
.dataB(s_logisimBus64[2:0]),
.result(s_logisimBus100[2:0]));
endmodule