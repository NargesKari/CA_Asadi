/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
mul11
**
**
**
*****************************************************************************/
module
mul11(
a,
b,
mul_out
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[31:0]
b;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[63:0]
mul_out;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus10;
wire
[63:0]
s_logisimBus100;
wire
[63:0]
s_logisimBus101;
wire
[63:0]
s_logisimBus102;
wire
[31:0]
s_logisimBus105;
wire
[63:0]
s_logisimBus106;
wire
[63:0]
s_logisimBus107;
wire
[63:0]
s_logisimBus108;
wire
[63:0]
s_logisimBus109;
wire
[31:0]
s_logisimBus110;
wire
[63:0]
s_logisimBus113;
wire
[63:0]
s_logisimBus114;
wire
[63:0]
s_logisimBus115;
wire
[63:0]
s_logisimBus116;
wire
[31:0]
s_logisimBus117;
wire
[31:0]
s_logisimBus120;
wire
[31:0]
s_logisimBus121;
wire
[63:0]
s_logisimBus122;
wire
[63:0]
s_logisimBus123;
wire
[63:0]
s_logisimBus124;
wire
[31:0]
s_logisimBus125;
wire
[31:0]
s_logisimBus128;
wire
[63:0]
s_logisimBus129;
wire
[31:0]
s_logisimBus13;
wire
[63:0]
s_logisimBus130;
wire
[63:0]
s_logisimBus131;
wire
[63:0]
s_logisimBus132;
wire
[63:0]
s_logisimBus135;
wire
[63:0]
s_logisimBus136;
wire
[31:0]
s_logisimBus137;
wire
[31:0]
s_logisimBus138;
wire
[31:0]
s_logisimBus139;
wire
[63:0]
s_logisimBus14;
wire
[63:0]
s_logisimBus140;
wire
[63:0]
s_logisimBus141;
wire
[31:0]
s_logisimBus142;
wire
[63:0]
s_logisimBus143;
wire
[63:0]
s_logisimBus144;
wire
[63:0]
s_logisimBus145;
wire
[63:0]
s_logisimBus146;
wire
[63:0]
s_logisimBus147;
wire
[63:0]
s_logisimBus148;
wire
[63:0]
s_logisimBus149;
wire
[31:0]
s_logisimBus15;
wire
[63:0]
s_logisimBus150;
wire
[63:0]
s_logisimBus151;
wire
[63:0]
s_logisimBus152;
wire
[63:0]
s_logisimBus153;
wire
[63:0]
s_logisimBus154;
wire
[63:0]
s_logisimBus155;
wire
[63:0]
s_logisimBus156;
wire
[63:0]
s_logisimBus157;
wire
[63:0]
s_logisimBus158;
wire
[63:0]
s_logisimBus159;
wire
[63:0]
s_logisimBus16;
wire
[63:0]
s_logisimBus160;
wire
[63:0]
s_logisimBus161;
wire
[63:0]
s_logisimBus162;
wire
[63:0]
s_logisimBus163;
wire
[63:0]
s_logisimBus164;
wire
[63:0]
s_logisimBus165;
wire
[63:0]
s_logisimBus166;
wire
[63:0]
s_logisimBus167;
wire
[63:0]
s_logisimBus168;
wire
[63:0]
s_logisimBus169;
wire
[63:0]
s_logisimBus17;
wire
[63:0]
s_logisimBus170;
wire
[63:0]
s_logisimBus171;
wire
[63:0]
s_logisimBus172;
wire
[63:0]
s_logisimBus173;
wire
[63:0]
s_logisimBus174;
wire
[63:0]
s_logisimBus175;
wire
[63:0]
s_logisimBus176;
wire
[63:0]
s_logisimBus177;
wire
[63:0]
s_logisimBus178;
wire
[63:0]
s_logisimBus179;
wire
[63:0]
s_logisimBus18;
wire
[31:0]
s_logisimBus180;
wire
[31:0]
s_logisimBus181;
wire
[63:0]
s_logisimBus19;
wire
[63:0]
s_logisimBus2;
wire
[63:0]
s_logisimBus20;
wire
[63:0]
s_logisimBus23;
wire
[63:0]
s_logisimBus24;
wire
[63:0]
s_logisimBus25;
wire
[63:0]
s_logisimBus26;
wire
[63:0]
s_logisimBus27;
wire
[63:0]
s_logisimBus28;
wire
[63:0]
s_logisimBus29;
wire
[31:0]
s_logisimBus3;
wire
[63:0]
s_logisimBus30;
wire
[63:0]
s_logisimBus31;
wire
[31:0]
s_logisimBus32;
wire
[31:0]
s_logisimBus35;
wire
[63:0]
s_logisimBus36;
wire
[63:0]
s_logisimBus37;
wire
[63:0]
s_logisimBus38;
wire
[63:0]
s_logisimBus39;
wire
[63:0]
s_logisimBus40;
wire
[31:0]
s_logisimBus41;
wire
[63:0]
s_logisimBus42;
wire
[63:0]
s_logisimBus45;
wire
[63:0]
s_logisimBus46;
wire
[63:0]
s_logisimBus47;
wire
[63:0]
s_logisimBus48;
wire
[31:0]
s_logisimBus49;
wire
[63:0]
s_logisimBus5;
wire
[31:0]
s_logisimBus52;
wire
[63:0]
s_logisimBus53;
wire
[63:0]
s_logisimBus54;
wire
[63:0]
s_logisimBus55;
wire
[63:0]
s_logisimBus56;
wire
[63:0]
s_logisimBus57;
wire
[63:0]
s_logisimBus58;
wire
[63:0]
s_logisimBus6;
wire
[31:0]
s_logisimBus61;
wire
[63:0]
s_logisimBus62;
wire
[63:0]
s_logisimBus63;
wire
[63:0]
s_logisimBus64;
wire
[63:0]
s_logisimBus65;
wire
[63:0]
s_logisimBus66;
wire
[63:0]
s_logisimBus67;
wire
[31:0]
s_logisimBus68;
wire
[63:0]
s_logisimBus7;
wire
[31:0]
s_logisimBus71;
wire
[63:0]
s_logisimBus72;
wire
[63:0]
s_logisimBus73;
wire
[63:0]
s_logisimBus74;
wire
[31:0]
s_logisimBus75;
wire
[31:0]
s_logisimBus76;
wire
[63:0]
s_logisimBus79;
wire
[31:0]
s_logisimBus8;
wire
[31:0]
s_logisimBus80;
wire
[63:0]
s_logisimBus81;
wire
[63:0]
s_logisimBus82;
wire
[63:0]
s_logisimBus83;
wire
[63:0]
s_logisimBus84;
wire
[63:0]
s_logisimBus87;
wire
[31:0]
s_logisimBus88;
wire
[63:0]
s_logisimBus89;
wire
[63:0]
s_logisimBus9;
wire
[63:0]
s_logisimBus90;
wire
[63:0]
s_logisimBus91;
wire
[63:0]
s_logisimBus92;
wire
[31:0]
s_logisimBus93;
wire
[31:0]
s_logisimBus94;
wire
[31:0]
s_logisimBus97;
wire
[63:0]
s_logisimBus98;
wire
[63:0]
s_logisimBus99;
wire
s_logisimNet1;
wire
s_logisimNet103;
wire
s_logisimNet104;
wire
s_logisimNet11;
wire
s_logisimNet111;
wire
s_logisimNet112;
wire
s_logisimNet118;
wire
s_logisimNet119;
wire
s_logisimNet12;
wire
s_logisimNet126;
wire
s_logisimNet127;
wire
s_logisimNet133;
wire
s_logisimNet134;
wire
s_logisimNet21;
wire
s_logisimNet22;
wire
s_logisimNet33;
wire
s_logisimNet34;
wire
s_logisimNet4;
wire
s_logisimNet43;
wire
s_logisimNet44;
wire
s_logisimNet50;
wire
s_logisimNet51;
wire
s_logisimNet59;
wire
s_logisimNet60;
wire
s_logisimNet69;
wire
s_logisimNet70;
wire
s_logisimNet77;
wire
s_logisimNet78;
wire
s_logisimNet85;
wire
s_logisimNet86;
wire
s_logisimNet95;
wire
s_logisimNet96;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus3[31:0]
=
a;
assign
s_logisimBus41[31:0]
=
b;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
mul_out
=
s_logisimBus113[63:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus25[63:0]
=
64'h0000000000000000;
assign
s_logisimBus65[63:0]
=
64'h0000000000000000;
assign
s_logisimBus24[63:0]
=
64'h0000000000000000;
assign
s_logisimBus52[31:0]
=
32'h00000013;
assign
s_logisimBus80[31:0]
=
32'h00000014;
assign
s_logisimBus105[31:0]
=
32'h00000015;
assign
s_logisimBus128[31:0]
=
32'h00000016;
assign
s_logisimBus0[31:0]
=
32'h00000017;
assign
s_logisimBus35[31:0]
=
32'h00000018;
assign
s_logisimBus71[31:0]
=
32'h00000019;
assign
s_logisimBus97[31:0]
=
32'h0000001A;
assign
s_logisimBus121[31:0]
=
32'h0000001B;
assign
s_logisimBus139[31:0]
=
32'h0000001C;
assign
s_logisimBus15[31:0]
=
32'h0000001D;
assign
s_logisimBus61[31:0]
=
32'h0000001E;
assign
s_logisimBus88[31:0]
=
32'h0000001F;
assign
s_logisimBus75[31:0]
=
32'h0000000E;
assign
s_logisimBus8[31:0]
=
32'h0000000A;
assign
s_logisimBus93[31:0]
=
32'h00000007;
assign
s_logisimBus137[31:0]
=
32'h00000009;
assign
s_logisimBus110[31:0]
=
32'h0000000B;
assign
s_logisimBus94[31:0]
=
32'h00000005;
assign
s_logisimBus117[31:0]
=
32'h00000006;
assign
s_logisimBus10[31:0]
=
32'h00000008;
assign
s_logisimBus49[31:0]
=
32'h0000000C;
assign
s_logisimBus76[31:0]
=
32'h0000000D;
assign
s_logisimBus125[31:0]
=
32'h0000000F;
assign
s_logisimBus142[31:0]
=
32'h00000010;
assign
s_logisimBus68[31:0]
=
32'h00000012;
assign
s_logisimBus32[31:0]
=
32'h00000001;
assign
s_logisimBus120[31:0]
=
32'h00000002;
assign
s_logisimBus138[31:0]
=
32'h00000003;
assign
s_logisimBus13[31:0]
=
32'h00000004;
assign
s_logisimBus180[31:0]
=
32'h00000011;
assign
s_logisimBus181[31:0]
=
32'h00000000;
assign
s_logisimBus148[63:0]
=
64'h0000000000000000;
assign
s_logisimBus149[63:0]
=
64'h0000000000000000;
assign
s_logisimBus150[63:0]
=
64'h0000000000000000;
assign
s_logisimBus151[63:0]
=
64'h0000000000000000;
assign
s_logisimBus152[63:0]
=
64'h0000000000000000;
assign
s_logisimBus153[63:0]
=
64'h0000000000000000;
assign
s_logisimBus154[63:0]
=
64'h0000000000000000;
assign
s_logisimBus155[63:0]
=
64'h0000000000000000;
assign
s_logisimBus156[63:0]
=
64'h0000000000000000;
assign
s_logisimBus157[63:0]
=
64'h0000000000000000;
assign
s_logisimBus158[63:0]
=
64'h0000000000000000;
assign
s_logisimBus159[63:0]
=
64'h0000000000000000;
assign
s_logisimBus160[63:0]
=
64'h0000000000000000;
assign
s_logisimBus161[63:0]
=
64'h0000000000000000;
assign
s_logisimBus162[63:0]
=
64'h0000000000000000;
assign
s_logisimBus163[63:0]
=
64'h0000000000000000;
assign
s_logisimBus164[63:0]
=
64'h0000000000000000;
assign
s_logisimBus165[63:0]
=
64'h0000000000000000;
assign
s_logisimBus166[63:0]
=
64'h0000000000000000;
assign
s_logisimBus167[63:0]
=
64'h0000000000000000;
assign
s_logisimBus168[63:0]
=
64'h0000000000000000;
assign
s_logisimBus169[63:0]
=
64'h0000000000000000;
assign
s_logisimBus170[63:0]
=
64'h0000000000000000;
assign
s_logisimBus171[63:0]
=
64'h0000000000000000;
assign
s_logisimBus172[63:0]
=
64'h0000000000000000;
assign
s_logisimBus173[63:0]
=
64'h0000000000000000;
assign
s_logisimBus174[63:0]
=
64'h0000000000000000;
assign
s_logisimBus175[63:0]
=
64'h0000000000000000;
assign
s_logisimBus176[63:0]
=
64'h0000000000000000;
assign
s_logisimBus177[63:0]
=
64'h0000000000000000;
assign
s_logisimBus178[63:0]
=
64'h0000000000000000;
assign
s_logisimBus179[63:0]
=
64'h0000000000000000;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_1
(.enable(1'b1),
.muxIn_0(s_logisimBus148[63:0]),
.muxIn_1(s_logisimBus36[63:0]),
.muxOut(s_logisimBus67[63:0]),
.sel(s_logisimBus41[10]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus149[63:0]),
.muxIn_1(s_logisimBus72[63:0]),
.muxOut(s_logisimBus19[63:0]),
.sel(s_logisimBus41[11]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus150[63:0]),
.muxIn_1(s_logisimBus98[63:0]),
.muxOut(s_logisimBus64[63:0]),
.sel(s_logisimBus41[12]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus151[63:0]),
.muxIn_1(s_logisimBus122[63:0]),
.muxOut(s_logisimBus91[63:0]),
.sel(s_logisimBus41[13]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus152[63:0]),
.muxIn_1(s_logisimBus140[63:0]),
.muxOut(s_logisimBus26[63:0]),
.sel(s_logisimBus41[14]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus153[63:0]),
.muxIn_1(s_logisimBus16[63:0]),
.muxOut(s_logisimBus6[63:0]),
.sel(s_logisimBus41[15]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_7
(.enable(1'b1),
.muxIn_0(s_logisimBus154[63:0]),
.muxIn_1(s_logisimBus62[63:0]),
.muxOut(s_logisimBus14[63:0]),
.sel(s_logisimBus41[16]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus155[63:0]),
.muxIn_1(s_logisimBus89[63:0]),
.muxOut(s_logisimBus79[63:0]),
.sel(s_logisimBus41[17]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_9
(.enable(1'b1),
.muxIn_0(s_logisimBus156[63:0]),
.muxIn_1(s_logisimBus114[63:0]),
.muxOut(s_logisimBus23[63:0]),
.sel(s_logisimBus41[18]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_10
(.enable(1'b1),
.muxIn_0(s_logisimBus157[63:0]),
.muxIn_1(s_logisimBus135[63:0]),
.muxOut(s_logisimBus92[63:0]),
.sel(s_logisimBus41[19]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_11
(.enable(1'b1),
.muxIn_0(s_logisimBus158[63:0]),
.muxIn_1(s_logisimBus146[63:0]),
.muxOut(s_logisimBus48[63:0]),
.sel(s_logisimBus41[20]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_12
(.enable(1'b1),
.muxIn_0(s_logisimBus159[63:0]),
.muxIn_1(s_logisimBus54[63:0]),
.muxOut(s_logisimBus20[63:0]),
.sel(s_logisimBus41[21]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_13
(.enable(1'b1),
.muxIn_0(s_logisimBus160[63:0]),
.muxIn_1(s_logisimBus82[63:0]),
.muxOut(s_logisimBus40[63:0]),
.sel(s_logisimBus41[22]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_14
(.enable(1'b1),
.muxIn_0(s_logisimBus161[63:0]),
.muxIn_1(s_logisimBus107[63:0]),
.muxOut(s_logisimBus74[63:0]),
.sel(s_logisimBus41[23]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_15
(.enable(1'b1),
.muxIn_0(s_logisimBus162[63:0]),
.muxIn_1(s_logisimBus130[63:0]),
.muxOut(s_logisimBus31[63:0]),
.sel(s_logisimBus41[24]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_16
(.enable(1'b1),
.muxIn_0(s_logisimBus163[63:0]),
.muxIn_1(s_logisimBus144[63:0]),
.muxOut(s_logisimBus57[63:0]),
.sel(s_logisimBus41[25]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_17
(.enable(1'b1),
.muxIn_0(s_logisimBus164[63:0]),
.muxIn_1(s_logisimBus37[63:0]),
.muxOut(s_logisimBus7[63:0]),
.sel(s_logisimBus41[26]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_18
(.enable(1'b1),
.muxIn_0(s_logisimBus165[63:0]),
.muxIn_1(s_logisimBus73[63:0]),
.muxOut(s_logisimBus5[63:0]),
.sel(s_logisimBus41[27]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_19
(.enable(1'b1),
.muxIn_0(s_logisimBus166[63:0]),
.muxIn_1(s_logisimBus99[63:0]),
.muxOut(s_logisimBus47[63:0]),
.sel(s_logisimBus41[28]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_20
(.enable(1'b1),
.muxIn_0(s_logisimBus167[63:0]),
.muxIn_1(s_logisimBus123[63:0]),
.muxOut(s_logisimBus56[63:0]),
.sel(s_logisimBus41[29]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_21
(.enable(1'b1),
.muxIn_0(s_logisimBus168[63:0]),
.muxIn_1(s_logisimBus141[63:0]),
.muxOut(s_logisimBus30[63:0]),
.sel(s_logisimBus41[30]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_22
(.enable(1'b1),
.muxIn_0(s_logisimBus169[63:0]),
.muxIn_1(s_logisimBus17[63:0]),
.muxOut(s_logisimBus9[63:0]),
.sel(s_logisimBus41[31]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_23
(.enable(1'b1),
.muxIn_0(s_logisimBus170[63:0]),
.muxIn_1(s_logisimBus63[63:0]),
.muxOut(s_logisimBus42[63:0]),
.sel(s_logisimBus41[0]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_24
(.enable(1'b1),
.muxIn_0(s_logisimBus171[63:0]),
.muxIn_1(s_logisimBus90[63:0]),
.muxOut(s_logisimBus55[63:0]),
.sel(s_logisimBus41[1]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_25
(.enable(1'b1),
.muxIn_0(s_logisimBus172[63:0]),
.muxIn_1(s_logisimBus115[63:0]),
.muxOut(s_logisimBus38[63:0]),
.sel(s_logisimBus41[2]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_26
(.enable(1'b1),
.muxIn_0(s_logisimBus173[63:0]),
.muxIn_1(s_logisimBus136[63:0]),
.muxOut(s_logisimBus108[63:0]),
.sel(s_logisimBus41[3]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_27
(.enable(1'b1),
.muxIn_0(s_logisimBus174[63:0]),
.muxIn_1(s_logisimBus147[63:0]),
.muxOut(s_logisimBus18[63:0]),
.sel(s_logisimBus41[4]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_28
(.enable(1'b1),
.muxIn_0(s_logisimBus175[63:0]),
.muxIn_1(s_logisimBus53[63:0]),
.muxOut(s_logisimBus29[63:0]),
.sel(s_logisimBus41[5]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_29
(.enable(1'b1),
.muxIn_0(s_logisimBus176[63:0]),
.muxIn_1(s_logisimBus81[63:0]),
.muxOut(s_logisimBus39[63:0]),
.sel(s_logisimBus41[6]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_30
(.enable(1'b1),
.muxIn_0(s_logisimBus177[63:0]),
.muxIn_1(s_logisimBus106[63:0]),
.muxOut(s_logisimBus2[63:0]),
.sel(s_logisimBus41[7]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_31
(.enable(1'b1),
.muxIn_0(s_logisimBus178[63:0]),
.muxIn_1(s_logisimBus129[63:0]),
.muxOut(s_logisimBus87[63:0]),
.sel(s_logisimBus41[8]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_32
(.enable(1'b1),
.muxIn_0(s_logisimBus179[63:0]),
.muxIn_1(s_logisimBus143[63:0]),
.muxOut(s_logisimBus27[63:0]),
.sel(s_logisimBus41[9]));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
CSaveA
CSaveA_15
(.a(s_logisimBus5[63:0]),
.b(s_logisimBus47[63:0]),
.c(s_logisimBus56[63:0]),
.sum(s_logisimBus58[63:0]));
CSaveA
CSaveA_17
(.a(s_logisimBus30[63:0]),
.b(s_logisimBus9[63:0]),
.c(s_logisimBus25[63:0]),
.sum(s_logisimBus83[63:0]));
CSaveA
CSaveA_5
(.a(s_logisimBus27[63:0]),
.b(s_logisimBus67[63:0]),
.c(s_logisimBus19[63:0]),
.sum(s_logisimBus132[63:0]));
CSaveA
CSaveA_9
(.a(s_logisimBus23[63:0]),
.b(s_logisimBus92[63:0]),
.c(s_logisimBus48[63:0]),
.sum(s_logisimBus45[63:0]));
CSaveA
CSaveA_12
(.a(s_logisimBus20[63:0]),
.b(s_logisimBus40[63:0]),
.c(s_logisimBus74[63:0]),
.sum(s_logisimBus66[63:0]));
CSaveA
CSaveA_1
(.a(s_logisimBus42[63:0]),
.b(s_logisimBus55[63:0]),
.c(s_logisimBus38[63:0]),
.sum(s_logisimBus84[63:0]));
CSaveA
CSaveA_3
(.a(s_logisimBus108[63:0]),
.b(s_logisimBus18[63:0]),
.c(s_logisimBus29[63:0]),
.sum(s_logisimBus102[63:0]));
CSaveA
CSaveA_4
(.a(s_logisimBus39[63:0]),
.b(s_logisimBus2[63:0]),
.c(s_logisimBus87[63:0]),
.sum(s_logisimBus46[63:0]));
CSaveA
CSaveA_7
(.a(s_logisimBus64[63:0]),
.b(s_logisimBus91[63:0]),
.c(s_logisimBus26[63:0]),
.sum(s_logisimBus28[63:0]));
CSaveA
CSaveA_13
(.a(s_logisimBus31[63:0]),
.b(s_logisimBus57[63:0]),
.c(s_logisimBus7[63:0]),
.sum(s_logisimBus131[63:0]));
CSaveA
CSaveA_8
(.a(s_logisimBus6[63:0]),
.b(s_logisimBus14[63:0]),
.c(s_logisimBus79[63:0]),
.sum(s_logisimBus100[63:0]));
CSaveA
CSaveA_6
(.a(s_logisimBus132[63:0]),
.b(s_logisimBus28[63:0]),
.c(s_logisimBus100[63:0]),
.sum(s_logisimBus124[63:0]));
CSaveA
CSaveA_11
(.a(s_logisimBus45[63:0]),
.b(s_logisimBus66[63:0]),
.c(s_logisimBus131[63:0]),
.sum(s_logisimBus109[63:0]));
CSaveA
CSaveA_16
(.a(s_logisimBus58[63:0]),
.b(s_logisimBus83[63:0]),
.c(s_logisimBus65[63:0]),
.sum(s_logisimBus116[63:0]));
CSaveA
CSaveA_2
(.a(s_logisimBus84[63:0]),
.b(s_logisimBus102[63:0]),
.c(s_logisimBus46[63:0]),
.sum(s_logisimBus101[63:0]));
CSaveA
CSaveA_10
(.a(s_logisimBus101[63:0]),
.b(s_logisimBus124[63:0]),
.c(s_logisimBus109[63:0]),
.sum(s_logisimBus145[63:0]));
CSaveA
CSaveA_14
(.a(s_logisimBus145[63:0]),
.b(s_logisimBus116[63:0]),
.c(s_logisimBus24[63:0]),
.sum(s_logisimBus113[63:0]));
SLL1
SLL1_11
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus8[31:0]),
.output1(s_logisimBus36[63:0]));
SLL1
SLL1_12
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus110[31:0]),
.output1(s_logisimBus72[63:0]));
SLL1
SLL1_13
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus49[31:0]),
.output1(s_logisimBus98[63:0]));
SLL1
SLL1_14
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus76[31:0]),
.output1(s_logisimBus122[63:0]));
SLL1
SLL1_15
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus75[31:0]),
.output1(s_logisimBus140[63:0]));
SLL1
SLL1_16
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus125[31:0]),
.output1(s_logisimBus16[63:0]));
SLL1
SLL1_17
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus142[31:0]),
.output1(s_logisimBus62[63:0]));
SLL1
SLL1_18
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus180[31:0]),
.output1(s_logisimBus89[63:0]));
SLL1
SLL1_19
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus68[31:0]),
.output1(s_logisimBus114[63:0]));
SLL1
SLL1_20
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus52[31:0]),
.output1(s_logisimBus135[63:0]));
SLL1
SLL1_21
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus80[31:0]),
.output1(s_logisimBus146[63:0]));
SLL1
SLL1_22
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus105[31:0]),
.output1(s_logisimBus54[63:0]));
SLL1
SLL1_23
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus128[31:0]),
.output1(s_logisimBus82[63:0]));
SLL1
SLL1_24
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus0[31:0]),
.output1(s_logisimBus107[63:0]));
SLL1
SLL1_25
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus35[31:0]),
.output1(s_logisimBus130[63:0]));
SLL1
SLL1_26
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus71[31:0]),
.output1(s_logisimBus144[63:0]));
SLL1
SLL1_27
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus97[31:0]),
.output1(s_logisimBus37[63:0]));
SLL1
SLL1_28
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus121[31:0]),
.output1(s_logisimBus73[63:0]));
SLL1
SLL1_29
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus139[31:0]),
.output1(s_logisimBus99[63:0]));
SLL1
SLL1_30
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus15[31:0]),
.output1(s_logisimBus123[63:0]));
SLL1
SLL1_31
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus61[31:0]),
.output1(s_logisimBus141[63:0]));
SLL1
SLL1_32
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus88[31:0]),
.output1(s_logisimBus17[63:0]));
SLL1
SLL1_1
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus181[31:0]),
.output1(s_logisimBus63[63:0]));
SLL1
SLL1_2
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus32[31:0]),
.output1(s_logisimBus90[63:0]));
SLL1
SLL1_3
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus120[31:0]),
.output1(s_logisimBus115[63:0]));
SLL1
SLL1_4
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus138[31:0]),
.output1(s_logisimBus136[63:0]));
SLL1
SLL1_5
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus13[31:0]),
.output1(s_logisimBus147[63:0]));
SLL1
SLL1_6
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus94[31:0]),
.output1(s_logisimBus53[63:0]));
SLL1
SLL1_7
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus117[31:0]),
.output1(s_logisimBus81[63:0]));
SLL1
SLL1_8
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus93[31:0]),
.output1(s_logisimBus106[63:0]));
SLL1
SLL1_9
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus10[31:0]),
.output1(s_logisimBus129[63:0]));
SLL1
SLL1_10
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus137[31:0]),
.output1(s_logisimBus143[63:0]));
endmodule