/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
inc_dec
**
**
**
*****************************************************************************/
module
inc_dec(
fuunc,
imm,
inc,
op,
rd,
rs,
rt,
shamt
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
inc;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[5:0]
fuunc;
output
[15:0]
imm;
output
[5:0]
op;
output
[4:0]
rd;
output
[4:0]
rs;
output
[4:0]
rt;
output
[4:0]
shamt;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[4:0]
s_logisimBus17;
wire
[4:0]
s_logisimBus18;
wire
[4:0]
s_logisimBus19;
wire
[5:0]
s_logisimBus23;
wire
[31:0]
s_logisimBus3;
wire
[4:0]
s_logisimBus35;
wire
[5:0]
s_logisimBus36;
wire
[15:0]
s_logisimBus37;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet10;
wire
s_logisimNet11;
wire
s_logisimNet12;
wire
s_logisimNet13;
wire
s_logisimNet14;
wire
s_logisimNet15;
wire
s_logisimNet16;
wire
s_logisimNet2;
wire
s_logisimNet20;
wire
s_logisimNet21;
wire
s_logisimNet22;
wire
s_logisimNet24;
wire
s_logisimNet25;
wire
s_logisimNet26;
wire
s_logisimNet27;
wire
s_logisimNet28;
wire
s_logisimNet29;
wire
s_logisimNet30;
wire
s_logisimNet31;
wire
s_logisimNet32;
wire
s_logisimNet33;
wire
s_logisimNet34;
wire
s_logisimNet38;
wire
s_logisimNet39;
wire
s_logisimNet4;
wire
s_logisimNet5;
wire
s_logisimNet6;
wire
s_logisimNet7;
wire
s_logisimNet8;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
wiring
is
defined
**
*******************************************************************************/
assign
s_logisimBus17[0]
=
s_logisimNet9;
assign
s_logisimBus17[1]
=
s_logisimNet26;
assign
s_logisimBus17[2]
=
s_logisimNet10;
assign
s_logisimBus17[3]
=
s_logisimNet27;
assign
s_logisimBus17[4]
=
s_logisimNet11;
assign
s_logisimBus18[0]
=
s_logisimNet20;
assign
s_logisimBus18[1]
=
s_logisimNet38;
assign
s_logisimBus18[2]
=
s_logisimNet21;
assign
s_logisimBus18[3]
=
s_logisimNet39;
assign
s_logisimBus18[4]
=
s_logisimNet22;
assign
s_logisimBus19[0]
=
s_logisimNet32;
assign
s_logisimBus19[1]
=
s_logisimNet15;
assign
s_logisimBus19[2]
=
s_logisimNet33;
assign
s_logisimBus19[3]
=
s_logisimNet16;
assign
s_logisimBus19[4]
=
s_logisimNet34;
assign
s_logisimBus23[0]
=
s_logisimNet25;
assign
s_logisimBus23[1]
=
s_logisimNet7;
assign
s_logisimBus23[2]
=
s_logisimNet24;
assign
s_logisimBus23[3]
=
s_logisimNet6;
assign
s_logisimBus23[4]
=
s_logisimNet28;
assign
s_logisimBus23[5]
=
s_logisimNet4;
assign
s_logisimBus35[0]
=
s_logisimNet0;
assign
s_logisimBus35[1]
=
s_logisimNet8;
assign
s_logisimBus35[2]
=
s_logisimNet1;
assign
s_logisimBus35[3]
=
s_logisimNet5;
assign
s_logisimBus35[4]
=
s_logisimNet2;
assign
s_logisimBus36[0]
=
s_logisimNet29;
assign
s_logisimBus36[1]
=
s_logisimNet12;
assign
s_logisimBus36[2]
=
s_logisimNet30;
assign
s_logisimBus36[3]
=
s_logisimNet13;
assign
s_logisimBus36[4]
=
s_logisimNet31;
assign
s_logisimBus36[5]
=
s_logisimNet14;
assign
s_logisimBus37[0]
=
s_logisimNet25;
assign
s_logisimBus37[10]
=
s_logisimNet2;
assign
s_logisimBus37[11]
=
s_logisimNet9;
assign
s_logisimBus37[12]
=
s_logisimNet26;
assign
s_logisimBus37[13]
=
s_logisimNet10;
assign
s_logisimBus37[14]
=
s_logisimNet27;
assign
s_logisimBus37[15]
=
s_logisimNet11;
assign
s_logisimBus37[1]
=
s_logisimNet7;
assign
s_logisimBus37[2]
=
s_logisimNet24;
assign
s_logisimBus37[3]
=
s_logisimNet6;
assign
s_logisimBus37[4]
=
s_logisimNet28;
assign
s_logisimBus37[5]
=
s_logisimNet4;
assign
s_logisimBus37[6]
=
s_logisimNet0;
assign
s_logisimBus37[7]
=
s_logisimNet8;
assign
s_logisimBus37[8]
=
s_logisimNet1;
assign
s_logisimBus37[9]
=
s_logisimNet5;
assign
s_logisimNet0
=
s_logisimBus3[6];
assign
s_logisimNet1
=
s_logisimBus3[8];
assign
s_logisimNet10
=
s_logisimBus3[13];
assign
s_logisimNet11
=
s_logisimBus3[15];
assign
s_logisimNet12
=
s_logisimBus3[27];
assign
s_logisimNet13
=
s_logisimBus3[29];
assign
s_logisimNet14
=
s_logisimBus3[31];
assign
s_logisimNet15
=
s_logisimBus3[22];
assign
s_logisimNet16
=
s_logisimBus3[24];
assign
s_logisimNet2
=
s_logisimBus3[10];
assign
s_logisimNet20
=
s_logisimBus3[16];
assign
s_logisimNet21
=
s_logisimBus3[18];
assign
s_logisimNet22
=
s_logisimBus3[20];
assign
s_logisimNet24
=
s_logisimBus3[2];
assign
s_logisimNet25
=
s_logisimBus3[0];
assign
s_logisimNet26
=
s_logisimBus3[12];
assign
s_logisimNet27
=
s_logisimBus3[14];
assign
s_logisimNet28
=
s_logisimBus3[4];
assign
s_logisimNet29
=
s_logisimBus3[26];
assign
s_logisimNet30
=
s_logisimBus3[28];
assign
s_logisimNet31
=
s_logisimBus3[30];
assign
s_logisimNet32
=
s_logisimBus3[21];
assign
s_logisimNet33
=
s_logisimBus3[23];
assign
s_logisimNet34
=
s_logisimBus3[25];
assign
s_logisimNet38
=
s_logisimBus3[17];
assign
s_logisimNet39
=
s_logisimBus3[19];
assign
s_logisimNet4
=
s_logisimBus3[5];
assign
s_logisimNet5
=
s_logisimBus3[9];
assign
s_logisimNet6
=
s_logisimBus3[3];
assign
s_logisimNet7
=
s_logisimBus3[1];
assign
s_logisimNet8
=
s_logisimBus3[7];
assign
s_logisimNet9
=
s_logisimBus3[11];
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus3[31:0]
=
inc;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
fuunc
=
s_logisimBus23[5:0];
assign
imm
=
s_logisimBus37[15:0];
assign
op
=
s_logisimBus36[5:0];
assign
rd
=
s_logisimBus17[4:0];
assign
rs
=
s_logisimBus19[4:0];
assign
rt
=
s_logisimBus18[4:0];
assign
shamt
=
s_logisimBus35[4:0];
endmodule