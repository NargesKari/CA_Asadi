/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
CU
**
**
**
*****************************************************************************/
module
CU(
ALUSrc,
AlUOp,
Branch,
IsNe,
Jump,
MemRead,
MemWrite,
MemtoReg,
RegDst,
RegWrite,
func,
isDiv,
isJal,
isMfhi,
isMflo,
isRJ,
isSll_shmt,
isSlti,
op_code
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[5:0]
func;
input
[5:0]
op_code;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
ALUSrc;
output
[3:0]
AlUOp;
output
Branch;
output
IsNe;
output
Jump;
output
MemRead;
output
MemWrite;
output
MemtoReg;
output
RegDst;
output
RegWrite;
output
isDiv;
output
isJal;
output
isMfhi;
output
isMflo;
output
isRJ;
output
isSll_shmt;
output
isSlti;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[3:0]
s_logisimBus60;
wire
[5:0]
s_logisimBus61;
wire
[5:0]
s_logisimBus62;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet10;
wire
s_logisimNet11;
wire
s_logisimNet12;
wire
s_logisimNet13;
wire
s_logisimNet14;
wire
s_logisimNet15;
wire
s_logisimNet16;
wire
s_logisimNet17;
wire
s_logisimNet18;
wire
s_logisimNet19;
wire
s_logisimNet2;
wire
s_logisimNet20;
wire
s_logisimNet21;
wire
s_logisimNet22;
wire
s_logisimNet23;
wire
s_logisimNet24;
wire
s_logisimNet25;
wire
s_logisimNet26;
wire
s_logisimNet27;
wire
s_logisimNet28;
wire
s_logisimNet29;
wire
s_logisimNet3;
wire
s_logisimNet30;
wire
s_logisimNet31;
wire
s_logisimNet32;
wire
s_logisimNet33;
wire
s_logisimNet34;
wire
s_logisimNet35;
wire
s_logisimNet36;
wire
s_logisimNet37;
wire
s_logisimNet38;
wire
s_logisimNet39;
wire
s_logisimNet4;
wire
s_logisimNet40;
wire
s_logisimNet41;
wire
s_logisimNet42;
wire
s_logisimNet43;
wire
s_logisimNet44;
wire
s_logisimNet45;
wire
s_logisimNet46;
wire
s_logisimNet47;
wire
s_logisimNet48;
wire
s_logisimNet49;
wire
s_logisimNet5;
wire
s_logisimNet50;
wire
s_logisimNet51;
wire
s_logisimNet52;
wire
s_logisimNet53;
wire
s_logisimNet54;
wire
s_logisimNet55;
wire
s_logisimNet56;
wire
s_logisimNet57;
wire
s_logisimNet58;
wire
s_logisimNet59;
wire
s_logisimNet6;
wire
s_logisimNet7;
wire
s_logisimNet8;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus61[5:0]
=
func;
assign
s_logisimBus62[5:0]
=
op_code;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
ALUSrc
=
s_logisimNet29;
assign
AlUOp
=
s_logisimBus60[3:0];
assign
Branch
=
s_logisimNet50;
assign
IsNe
=
s_logisimNet40;
assign
Jump
=
s_logisimNet44;
assign
MemRead
=
s_logisimNet7;
assign
MemWrite
=
s_logisimNet28;
assign
MemtoReg
=
s_logisimNet7;
assign
RegDst
=
s_logisimNet35;
assign
RegWrite
=
s_logisimNet8;
assign
isDiv
=
s_logisimNet47;
assign
isJal
=
s_logisimNet24;
assign
isMfhi
=
s_logisimNet4;
assign
isMflo
=
s_logisimNet39;
assign
isRJ
=
s_logisimNet53;
assign
isSll_shmt
=
s_logisimNet36;
assign
isSlti
=
s_logisimNet32;
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimNet19
=
~s_logisimBus61[5];
assign
s_logisimNet9
=
~s_logisimBus61[4];
assign
s_logisimNet17
=
~s_logisimBus61[3];
assign
s_logisimNet13
=
~s_logisimBus61[2];
assign
s_logisimNet26
=
~s_logisimBus61[1];
assign
s_logisimNet10
=
~s_logisimBus61[0];
assign
s_logisimNet6
=
~s_logisimBus62[5];
assign
s_logisimNet15
=
~s_logisimBus62[4];
assign
s_logisimNet31
=
~s_logisimBus62[3];
assign
s_logisimNet27
=
~s_logisimBus62[2];
assign
s_logisimNet11
=
~s_logisimBus62[1];
assign
s_logisimNet0
=
~s_logisimBus62[0];
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE_5_INPUTS
#(.BubblesMask({1'b0,
4'h0}))
GATES_1
(.input1(s_logisimNet28),
.input2(s_logisimNet25),
.input3(1'b0),
.input4(s_logisimNet7),
.input5(s_logisimNet32),
.result(s_logisimNet29));
OR_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
GATES_2
(.input1(s_logisimNet3),
.input2(s_logisimNet7),
.input3(s_logisimNet34),
.input4(s_logisimNet25),
.input5(s_logisimNet32),
.input6(s_logisimNet24),
.result(s_logisimNet46));
AND_GATE
#(.BubblesMask(2'b00))
GATES_3
(.input1(s_logisimNet46),
.input2(s_logisimNet38),
.result(s_logisimNet8));
NOR_GATE
#(.BubblesMask(2'b00))
GATES_4
(.input1(s_logisimNet47),
.input2(s_logisimNet53),
.result(s_logisimNet38));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
mfloo
(.input1(s_logisimNet3),
.input2(s_logisimNet10),
.input3(s_logisimBus61[1]),
.input4(s_logisimNet13),
.input5(s_logisimNet17),
.input6(s_logisimBus61[4]),
.input7(s_logisimNet19),
.result(s_logisimNet39));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
div
(.input1(s_logisimNet3),
.input2(s_logisimNet10),
.input3(s_logisimBus61[1]),
.input4(s_logisimNet13),
.input5(s_logisimBus61[3]),
.input6(s_logisimBus61[4]),
.input7(s_logisimNet19),
.result(s_logisimNet47));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
sll_old
(.input1(s_logisimNet3),
.input2(s_logisimNet10),
.input3(s_logisimNet26),
.input4(s_logisimBus61[2]),
.input5(s_logisimNet17),
.input6(s_logisimNet9),
.input7(s_logisimNet19),
.result(s_logisimNet57));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
jr
(.input1(s_logisimNet3),
.input2(s_logisimNet10),
.input3(s_logisimNet26),
.input4(s_logisimNet13),
.input5(s_logisimBus61[3]),
.input6(s_logisimNet9),
.input7(s_logisimNet19),
.result(s_logisimNet53));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
mul
(.input1(s_logisimNet34),
.input2(s_logisimNet10),
.input3(s_logisimBus61[1]),
.input4(s_logisimNet13),
.input5(s_logisimNet17),
.input6(s_logisimNet9),
.input7(s_logisimNet19),
.result(s_logisimNet49));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
add
(.input1(s_logisimNet3),
.input2(s_logisimNet10),
.input3(s_logisimNet26),
.input4(s_logisimNet13),
.input5(s_logisimNet17),
.input6(s_logisimNet9),
.input7(s_logisimBus61[5]),
.result(s_logisimNet45));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
sub
(.input1(s_logisimNet3),
.input2(s_logisimNet10),
.input3(s_logisimBus61[1]),
.input4(s_logisimNet13),
.input5(s_logisimNet17),
.input6(s_logisimNet9),
.input7(s_logisimBus61[5]),
.result(s_logisimNet18));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
annd
(.input1(s_logisimNet3),
.input2(s_logisimNet10),
.input3(s_logisimNet26),
.input4(s_logisimBus61[2]),
.input5(s_logisimNet17),
.input6(s_logisimNet9),
.input7(s_logisimBus61[5]),
.result(s_logisimNet56));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
Or1
(.input1(s_logisimNet3),
.input2(s_logisimBus61[0]),
.input3(s_logisimNet26),
.input4(s_logisimBus61[2]),
.input5(s_logisimNet17),
.input6(s_logisimNet9),
.input7(s_logisimBus61[5]),
.result(s_logisimNet54));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
xor1
(.input1(s_logisimNet3),
.input2(s_logisimNet10),
.input3(s_logisimBus61[1]),
.input4(s_logisimBus61[2]),
.input5(s_logisimNet17),
.input6(s_logisimNet9),
.input7(s_logisimBus61[5]),
.result(s_logisimNet58));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
sll_SH
(.input1(s_logisimNet3),
.input2(s_logisimNet10),
.input3(s_logisimNet26),
.input4(s_logisimNet13),
.input5(s_logisimNet17),
.input6(s_logisimNet9),
.input7(s_logisimNet19),
.result(s_logisimNet36));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
srl1
(.input1(s_logisimNet3),
.input2(s_logisimNet10),
.input3(s_logisimBus61[1]),
.input4(s_logisimBus61[2]),
.input5(s_logisimNet17),
.input6(s_logisimNet9),
.input7(s_logisimNet19),
.result(s_logisimNet52));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
sra1
(.input1(s_logisimNet3),
.input2(s_logisimBus61[0]),
.input3(s_logisimBus61[1]),
.input4(s_logisimBus61[2]),
.input5(s_logisimNet17),
.input6(s_logisimNet9),
.input7(s_logisimNet19),
.result(s_logisimNet59));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
mfhii
(.input1(s_logisimNet3),
.input2(s_logisimNet10),
.input3(s_logisimNet26),
.input4(s_logisimNet13),
.input5(s_logisimNet17),
.input6(s_logisimBus61[4]),
.input7(s_logisimNet19),
.result(s_logisimNet4));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
jal
(.input1(s_logisimNet6),
.input2(s_logisimNet15),
.input3(s_logisimNet31),
.input4(s_logisimNet27),
.input5(s_logisimBus62[1]),
.input6(s_logisimBus62[0]),
.result(s_logisimNet24));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
beq
(.input1(s_logisimNet6),
.input2(s_logisimNet15),
.input3(s_logisimNet31),
.input4(s_logisimBus62[2]),
.input5(s_logisimNet11),
.input6(s_logisimNet0),
.result(s_logisimNet51));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
R_type
(.input1(s_logisimNet0),
.input2(s_logisimNet11),
.input3(s_logisimNet27),
.input4(s_logisimNet31),
.input5(s_logisimNet15),
.input6(s_logisimNet6),
.result(s_logisimNet3));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
addi
(.input1(s_logisimNet0),
.input2(s_logisimNet11),
.input3(s_logisimNet27),
.input4(s_logisimBus62[3]),
.input5(s_logisimNet15),
.input6(s_logisimNet6),
.result(s_logisimNet25));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
sw
(.input1(s_logisimBus62[0]),
.input2(s_logisimBus62[1]),
.input3(s_logisimNet27),
.input4(s_logisimBus62[3]),
.input5(s_logisimNet15),
.input6(s_logisimBus62[5]),
.result(s_logisimNet28));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
lw
(.input1(s_logisimBus62[5]),
.input2(s_logisimNet15),
.input3(s_logisimNet31),
.input4(s_logisimNet27),
.input5(s_logisimBus62[1]),
.input6(s_logisimBus62[0]),
.result(s_logisimNet7));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
bne
(.input1(s_logisimNet6),
.input2(s_logisimNet15),
.input3(s_logisimNet31),
.input4(s_logisimBus62[2]),
.input5(s_logisimNet11),
.input6(s_logisimBus62[0]),
.result(s_logisimNet40));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
slti
(.input1(s_logisimNet6),
.input2(s_logisimNet15),
.input3(s_logisimBus62[3]),
.input4(s_logisimNet27),
.input5(s_logisimBus62[1]),
.input6(s_logisimNet0),
.result(s_logisimNet32));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
j
(.input1(s_logisimNet6),
.input2(s_logisimNet15),
.input3(s_logisimNet31),
.input4(s_logisimNet27),
.input5(s_logisimBus62[1]),
.input6(s_logisimNet0),
.result(s_logisimNet21));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
mul1
(.input1(s_logisimNet6),
.input2(s_logisimBus62[4]),
.input3(s_logisimBus62[3]),
.input4(s_logisimBus62[2]),
.input5(s_logisimNet11),
.input6(s_logisimNet0),
.result(s_logisimNet34));
OR_GATE
#(.BubblesMask(2'b00))
GATES_29
(.input1(s_logisimNet3),
.input2(s_logisimNet34),
.result(s_logisimNet35));
OR_GATE_3_INPUTS
#(.BubblesMask(3'b000))
GATES_30
(.input1(s_logisimNet21),
.input2(s_logisimNet24),
.input3(s_logisimNet53),
.result(s_logisimNet44));
OR_GATE
#(.BubblesMask(2'b00))
GATES_31
(.input1(s_logisimNet40),
.input2(s_logisimNet51),
.result(s_logisimNet42));
OR_GATE
#(.BubblesMask(2'b00))
GATES_32
(.input1(s_logisimNet40),
.input2(s_logisimNet51),
.result(s_logisimNet50));
OR_GATE_5_INPUTS
#(.BubblesMask({1'b0,
4'h0}))
GATES_33
(.input1(s_logisimNet52),
.input2(s_logisimNet59),
.input3(s_logisimNet49),
.input4(s_logisimNet47),
.input5(s_logisimNet58),
.result(s_logisimBus60[1]));
OR_GATE_3_INPUTS
#(.BubblesMask(3'b000))
GATES_34
(.input1(s_logisimNet56),
.input2(s_logisimNet54),
.input3(s_logisimNet58),
.result(s_logisimBus60[2]));
OR_GATE_4_INPUTS
#(.BubblesMask(4'h0))
GATES_35
(.input1(s_logisimNet57),
.input2(s_logisimNet59),
.input3(s_logisimNet52),
.input4(s_logisimNet36),
.result(s_logisimBus60[3]));
OR_GATE_8_INPUTS
#(.BubblesMask(8'h00))
GATES_36
(.input1(s_logisimNet54),
.input2(s_logisimNet42),
.input3(s_logisimNet47),
.input4(s_logisimNet18),
.input5(s_logisimNet36),
.input6(s_logisimNet59),
.input7(s_logisimNet57),
.input8(s_logisimNet32),
.result(s_logisimBus60[0]));
endmodule