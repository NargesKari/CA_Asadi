/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
ALU_CSA
**
**
**
*****************************************************************************/
module
ALU_CSA(
A,
B,
SUM,
cin,
cout
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
A;
input
[31:0]
B;
input
cin;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[31:0]
SUM;
output
cout;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[7:0]
s_logisimBus11;
wire
[7:0]
s_logisimBus20;
wire
[7:0]
s_logisimBus23;
wire
[7:0]
s_logisimBus24;
wire
[7:0]
s_logisimBus26;
wire
[31:0]
s_logisimBus27;
wire
[31:0]
s_logisimBus31;
wire
[31:0]
s_logisimBus32;
wire
[7:0]
s_logisimBus7;
wire
s_logisimNet10;
wire
s_logisimNet12;
wire
s_logisimNet16;
wire
s_logisimNet19;
wire
s_logisimNet2;
wire
s_logisimNet28;
wire
s_logisimNet29;
wire
s_logisimNet3;
wire
s_logisimNet30;
wire
s_logisimNet4;
wire
s_logisimNet5;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus31[31:0]
=
A;
assign
s_logisimBus32[31:0]
=
B;
assign
s_logisimNet3
=
cin;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
SUM
=
s_logisimBus27[31:0];
assign
cout
=
s_logisimNet28;
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimNet4
=
1'b1;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Multiplexer_bus_2
#(.nrOfBits(8))
PLEXERS_1
(.enable(1'b1),
.muxIn_0(s_logisimBus23[7:0]),
.muxIn_1(s_logisimBus24[7:0]),
.muxOut(s_logisimBus27[15:8]),
.sel(s_logisimNet9));
Multiplexer_2
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimNet16),
.muxIn_1(s_logisimNet2),
.muxOut(s_logisimNet12),
.sel(s_logisimNet9));
Multiplexer_bus_2
#(.nrOfBits(8))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus7[7:0]),
.muxIn_1(s_logisimBus11[7:0]),
.muxOut(s_logisimBus27[23:16]),
.sel(s_logisimNet12));
Multiplexer_2
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimNet30),
.muxIn_1(s_logisimNet5),
.muxOut(s_logisimNet10),
.sel(s_logisimNet12));
Multiplexer_bus_2
#(.nrOfBits(8))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus26[7:0]),
.muxIn_1(s_logisimBus20[7:0]),
.muxOut(s_logisimBus27[31:24]),
.sel(s_logisimNet10));
Multiplexer_2
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimNet19),
.muxIn_1(s_logisimNet29),
.muxOut(s_logisimNet28),
.sel(s_logisimNet10));
Adder
#(.extendedBits(9),
.nrOfBits(8))
ARITH_7
(.carryIn(s_logisimNet3),
.carryOut(s_logisimNet9),
.dataA(s_logisimBus31[7:0]),
.dataB(s_logisimBus32[7:0]),
.result(s_logisimBus27[7:0]));
Adder
#(.extendedBits(9),
.nrOfBits(8))
ARITH_8
(.carryIn(1'b0),
.carryOut(s_logisimNet30),
.dataA(s_logisimBus31[23:16]),
.dataB(s_logisimBus32[23:16]),
.result(s_logisimBus7[7:0]));
Adder
#(.extendedBits(9),
.nrOfBits(8))
ARITH_9
(.carryIn(1'b0),
.carryOut(s_logisimNet16),
.dataA(s_logisimBus31[15:8]),
.dataB(s_logisimBus32[15:8]),
.result(s_logisimBus23[7:0]));
Adder
#(.extendedBits(9),
.nrOfBits(8))
ARITH_10
(.carryIn(s_logisimNet4),
.carryOut(s_logisimNet2),
.dataA(s_logisimBus31[15:8]),
.dataB(s_logisimBus32[15:8]),
.result(s_logisimBus24[7:0]));
Adder
#(.extendedBits(9),
.nrOfBits(8))
ARITH_11
(.carryIn(s_logisimNet4),
.carryOut(s_logisimNet5),
.dataA(s_logisimBus31[23:16]),
.dataB(s_logisimBus32[23:16]),
.result(s_logisimBus11[7:0]));
Adder
#(.extendedBits(9),
.nrOfBits(8))
ARITH_12
(.carryIn(1'b0),
.carryOut(s_logisimNet19),
.dataA(s_logisimBus31[31:24]),
.dataB(s_logisimBus32[31:24]),
.result(s_logisimBus26[7:0]));
Adder
#(.extendedBits(9),
.nrOfBits(8))
ARITH_13
(.carryIn(s_logisimNet4),
.carryOut(s_logisimNet29),
.dataA(s_logisimBus31[31:24]),
.dataB(s_logisimBus32[31:24]),
.result(s_logisimBus20[7:0]));
endmodule