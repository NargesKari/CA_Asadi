/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
ALU_CSaveA
**
**
**
*****************************************************************************/
module
ALU_CSaveA(
a,
b,
c,
sum
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[63:0]
a;
input
[63:0]
b;
input
[63:0]
c;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[63:0]
sum;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[63:0]
s_logisimBus227;
wire
[63:0]
s_logisimBus283;
wire
[63:0]
s_logisimBus443;
wire
[63:0]
s_logisimBus448;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet10;
wire
s_logisimNet100;
wire
s_logisimNet101;
wire
s_logisimNet102;
wire
s_logisimNet103;
wire
s_logisimNet104;
wire
s_logisimNet105;
wire
s_logisimNet106;
wire
s_logisimNet107;
wire
s_logisimNet108;
wire
s_logisimNet109;
wire
s_logisimNet11;
wire
s_logisimNet110;
wire
s_logisimNet111;
wire
s_logisimNet112;
wire
s_logisimNet113;
wire
s_logisimNet114;
wire
s_logisimNet115;
wire
s_logisimNet116;
wire
s_logisimNet117;
wire
s_logisimNet118;
wire
s_logisimNet119;
wire
s_logisimNet12;
wire
s_logisimNet120;
wire
s_logisimNet121;
wire
s_logisimNet122;
wire
s_logisimNet123;
wire
s_logisimNet124;
wire
s_logisimNet125;
wire
s_logisimNet126;
wire
s_logisimNet127;
wire
s_logisimNet128;
wire
s_logisimNet129;
wire
s_logisimNet13;
wire
s_logisimNet130;
wire
s_logisimNet131;
wire
s_logisimNet132;
wire
s_logisimNet133;
wire
s_logisimNet134;
wire
s_logisimNet135;
wire
s_logisimNet136;
wire
s_logisimNet137;
wire
s_logisimNet138;
wire
s_logisimNet139;
wire
s_logisimNet14;
wire
s_logisimNet140;
wire
s_logisimNet141;
wire
s_logisimNet142;
wire
s_logisimNet143;
wire
s_logisimNet144;
wire
s_logisimNet145;
wire
s_logisimNet146;
wire
s_logisimNet147;
wire
s_logisimNet148;
wire
s_logisimNet149;
wire
s_logisimNet15;
wire
s_logisimNet150;
wire
s_logisimNet151;
wire
s_logisimNet152;
wire
s_logisimNet153;
wire
s_logisimNet154;
wire
s_logisimNet155;
wire
s_logisimNet156;
wire
s_logisimNet157;
wire
s_logisimNet158;
wire
s_logisimNet159;
wire
s_logisimNet16;
wire
s_logisimNet160;
wire
s_logisimNet161;
wire
s_logisimNet162;
wire
s_logisimNet163;
wire
s_logisimNet164;
wire
s_logisimNet165;
wire
s_logisimNet166;
wire
s_logisimNet167;
wire
s_logisimNet168;
wire
s_logisimNet169;
wire
s_logisimNet17;
wire
s_logisimNet170;
wire
s_logisimNet171;
wire
s_logisimNet172;
wire
s_logisimNet173;
wire
s_logisimNet174;
wire
s_logisimNet175;
wire
s_logisimNet176;
wire
s_logisimNet177;
wire
s_logisimNet178;
wire
s_logisimNet179;
wire
s_logisimNet18;
wire
s_logisimNet180;
wire
s_logisimNet181;
wire
s_logisimNet182;
wire
s_logisimNet183;
wire
s_logisimNet184;
wire
s_logisimNet185;
wire
s_logisimNet186;
wire
s_logisimNet187;
wire
s_logisimNet188;
wire
s_logisimNet189;
wire
s_logisimNet19;
wire
s_logisimNet190;
wire
s_logisimNet191;
wire
s_logisimNet192;
wire
s_logisimNet193;
wire
s_logisimNet194;
wire
s_logisimNet195;
wire
s_logisimNet196;
wire
s_logisimNet197;
wire
s_logisimNet198;
wire
s_logisimNet199;
wire
s_logisimNet2;
wire
s_logisimNet20;
wire
s_logisimNet200;
wire
s_logisimNet201;
wire
s_logisimNet202;
wire
s_logisimNet203;
wire
s_logisimNet204;
wire
s_logisimNet205;
wire
s_logisimNet206;
wire
s_logisimNet207;
wire
s_logisimNet208;
wire
s_logisimNet209;
wire
s_logisimNet21;
wire
s_logisimNet210;
wire
s_logisimNet211;
wire
s_logisimNet212;
wire
s_logisimNet213;
wire
s_logisimNet214;
wire
s_logisimNet215;
wire
s_logisimNet216;
wire
s_logisimNet217;
wire
s_logisimNet218;
wire
s_logisimNet219;
wire
s_logisimNet22;
wire
s_logisimNet220;
wire
s_logisimNet221;
wire
s_logisimNet222;
wire
s_logisimNet223;
wire
s_logisimNet224;
wire
s_logisimNet225;
wire
s_logisimNet226;
wire
s_logisimNet228;
wire
s_logisimNet229;
wire
s_logisimNet23;
wire
s_logisimNet230;
wire
s_logisimNet231;
wire
s_logisimNet232;
wire
s_logisimNet233;
wire
s_logisimNet234;
wire
s_logisimNet235;
wire
s_logisimNet236;
wire
s_logisimNet237;
wire
s_logisimNet238;
wire
s_logisimNet239;
wire
s_logisimNet24;
wire
s_logisimNet240;
wire
s_logisimNet241;
wire
s_logisimNet242;
wire
s_logisimNet243;
wire
s_logisimNet244;
wire
s_logisimNet245;
wire
s_logisimNet246;
wire
s_logisimNet247;
wire
s_logisimNet248;
wire
s_logisimNet249;
wire
s_logisimNet25;
wire
s_logisimNet250;
wire
s_logisimNet251;
wire
s_logisimNet252;
wire
s_logisimNet253;
wire
s_logisimNet254;
wire
s_logisimNet255;
wire
s_logisimNet256;
wire
s_logisimNet257;
wire
s_logisimNet258;
wire
s_logisimNet259;
wire
s_logisimNet26;
wire
s_logisimNet260;
wire
s_logisimNet261;
wire
s_logisimNet262;
wire
s_logisimNet263;
wire
s_logisimNet264;
wire
s_logisimNet265;
wire
s_logisimNet266;
wire
s_logisimNet267;
wire
s_logisimNet268;
wire
s_logisimNet269;
wire
s_logisimNet27;
wire
s_logisimNet270;
wire
s_logisimNet271;
wire
s_logisimNet272;
wire
s_logisimNet273;
wire
s_logisimNet274;
wire
s_logisimNet275;
wire
s_logisimNet276;
wire
s_logisimNet277;
wire
s_logisimNet278;
wire
s_logisimNet279;
wire
s_logisimNet28;
wire
s_logisimNet280;
wire
s_logisimNet281;
wire
s_logisimNet282;
wire
s_logisimNet284;
wire
s_logisimNet285;
wire
s_logisimNet286;
wire
s_logisimNet287;
wire
s_logisimNet288;
wire
s_logisimNet289;
wire
s_logisimNet29;
wire
s_logisimNet290;
wire
s_logisimNet291;
wire
s_logisimNet292;
wire
s_logisimNet293;
wire
s_logisimNet294;
wire
s_logisimNet295;
wire
s_logisimNet296;
wire
s_logisimNet297;
wire
s_logisimNet298;
wire
s_logisimNet299;
wire
s_logisimNet3;
wire
s_logisimNet30;
wire
s_logisimNet300;
wire
s_logisimNet301;
wire
s_logisimNet302;
wire
s_logisimNet303;
wire
s_logisimNet304;
wire
s_logisimNet305;
wire
s_logisimNet306;
wire
s_logisimNet307;
wire
s_logisimNet308;
wire
s_logisimNet309;
wire
s_logisimNet31;
wire
s_logisimNet310;
wire
s_logisimNet311;
wire
s_logisimNet312;
wire
s_logisimNet313;
wire
s_logisimNet314;
wire
s_logisimNet315;
wire
s_logisimNet316;
wire
s_logisimNet317;
wire
s_logisimNet318;
wire
s_logisimNet319;
wire
s_logisimNet32;
wire
s_logisimNet320;
wire
s_logisimNet321;
wire
s_logisimNet322;
wire
s_logisimNet323;
wire
s_logisimNet324;
wire
s_logisimNet325;
wire
s_logisimNet326;
wire
s_logisimNet327;
wire
s_logisimNet328;
wire
s_logisimNet329;
wire
s_logisimNet33;
wire
s_logisimNet330;
wire
s_logisimNet331;
wire
s_logisimNet332;
wire
s_logisimNet333;
wire
s_logisimNet334;
wire
s_logisimNet335;
wire
s_logisimNet336;
wire
s_logisimNet337;
wire
s_logisimNet338;
wire
s_logisimNet339;
wire
s_logisimNet34;
wire
s_logisimNet340;
wire
s_logisimNet341;
wire
s_logisimNet342;
wire
s_logisimNet343;
wire
s_logisimNet344;
wire
s_logisimNet345;
wire
s_logisimNet346;
wire
s_logisimNet347;
wire
s_logisimNet348;
wire
s_logisimNet349;
wire
s_logisimNet35;
wire
s_logisimNet350;
wire
s_logisimNet351;
wire
s_logisimNet352;
wire
s_logisimNet353;
wire
s_logisimNet354;
wire
s_logisimNet355;
wire
s_logisimNet356;
wire
s_logisimNet357;
wire
s_logisimNet358;
wire
s_logisimNet359;
wire
s_logisimNet36;
wire
s_logisimNet360;
wire
s_logisimNet361;
wire
s_logisimNet362;
wire
s_logisimNet363;
wire
s_logisimNet364;
wire
s_logisimNet365;
wire
s_logisimNet366;
wire
s_logisimNet367;
wire
s_logisimNet368;
wire
s_logisimNet369;
wire
s_logisimNet37;
wire
s_logisimNet370;
wire
s_logisimNet371;
wire
s_logisimNet372;
wire
s_logisimNet373;
wire
s_logisimNet374;
wire
s_logisimNet375;
wire
s_logisimNet376;
wire
s_logisimNet377;
wire
s_logisimNet378;
wire
s_logisimNet379;
wire
s_logisimNet38;
wire
s_logisimNet380;
wire
s_logisimNet381;
wire
s_logisimNet382;
wire
s_logisimNet383;
wire
s_logisimNet384;
wire
s_logisimNet385;
wire
s_logisimNet386;
wire
s_logisimNet387;
wire
s_logisimNet388;
wire
s_logisimNet389;
wire
s_logisimNet39;
wire
s_logisimNet390;
wire
s_logisimNet391;
wire
s_logisimNet392;
wire
s_logisimNet393;
wire
s_logisimNet394;
wire
s_logisimNet395;
wire
s_logisimNet396;
wire
s_logisimNet397;
wire
s_logisimNet398;
wire
s_logisimNet399;
wire
s_logisimNet4;
wire
s_logisimNet40;
wire
s_logisimNet400;
wire
s_logisimNet401;
wire
s_logisimNet402;
wire
s_logisimNet403;
wire
s_logisimNet404;
wire
s_logisimNet405;
wire
s_logisimNet406;
wire
s_logisimNet407;
wire
s_logisimNet408;
wire
s_logisimNet409;
wire
s_logisimNet41;
wire
s_logisimNet410;
wire
s_logisimNet411;
wire
s_logisimNet412;
wire
s_logisimNet413;
wire
s_logisimNet414;
wire
s_logisimNet415;
wire
s_logisimNet416;
wire
s_logisimNet417;
wire
s_logisimNet418;
wire
s_logisimNet419;
wire
s_logisimNet42;
wire
s_logisimNet420;
wire
s_logisimNet421;
wire
s_logisimNet422;
wire
s_logisimNet423;
wire
s_logisimNet424;
wire
s_logisimNet425;
wire
s_logisimNet426;
wire
s_logisimNet427;
wire
s_logisimNet428;
wire
s_logisimNet429;
wire
s_logisimNet43;
wire
s_logisimNet430;
wire
s_logisimNet431;
wire
s_logisimNet432;
wire
s_logisimNet433;
wire
s_logisimNet434;
wire
s_logisimNet435;
wire
s_logisimNet436;
wire
s_logisimNet437;
wire
s_logisimNet438;
wire
s_logisimNet439;
wire
s_logisimNet44;
wire
s_logisimNet440;
wire
s_logisimNet441;
wire
s_logisimNet442;
wire
s_logisimNet444;
wire
s_logisimNet445;
wire
s_logisimNet446;
wire
s_logisimNet447;
wire
s_logisimNet45;
wire
s_logisimNet46;
wire
s_logisimNet47;
wire
s_logisimNet48;
wire
s_logisimNet49;
wire
s_logisimNet5;
wire
s_logisimNet50;
wire
s_logisimNet51;
wire
s_logisimNet52;
wire
s_logisimNet53;
wire
s_logisimNet54;
wire
s_logisimNet55;
wire
s_logisimNet56;
wire
s_logisimNet57;
wire
s_logisimNet58;
wire
s_logisimNet59;
wire
s_logisimNet6;
wire
s_logisimNet60;
wire
s_logisimNet61;
wire
s_logisimNet62;
wire
s_logisimNet63;
wire
s_logisimNet64;
wire
s_logisimNet65;
wire
s_logisimNet66;
wire
s_logisimNet67;
wire
s_logisimNet68;
wire
s_logisimNet69;
wire
s_logisimNet7;
wire
s_logisimNet70;
wire
s_logisimNet71;
wire
s_logisimNet72;
wire
s_logisimNet73;
wire
s_logisimNet74;
wire
s_logisimNet75;
wire
s_logisimNet76;
wire
s_logisimNet77;
wire
s_logisimNet78;
wire
s_logisimNet79;
wire
s_logisimNet8;
wire
s_logisimNet80;
wire
s_logisimNet81;
wire
s_logisimNet82;
wire
s_logisimNet83;
wire
s_logisimNet84;
wire
s_logisimNet85;
wire
s_logisimNet86;
wire
s_logisimNet87;
wire
s_logisimNet88;
wire
s_logisimNet89;
wire
s_logisimNet9;
wire
s_logisimNet90;
wire
s_logisimNet91;
wire
s_logisimNet92;
wire
s_logisimNet93;
wire
s_logisimNet94;
wire
s_logisimNet95;
wire
s_logisimNet96;
wire
s_logisimNet97;
wire
s_logisimNet98;
wire
s_logisimNet99;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus227[63:0]
=
b;
assign
s_logisimBus283[63:0]
=
c;
assign
s_logisimBus443[63:0]
=
a;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
sum
=
s_logisimBus448[63:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimNet444
=
1'b0;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
FullAdder
#(.extendedBits(2))
ARITH_1
(.carryIn(s_logisimBus443[10]),
.carryOut(s_logisimNet79),
.dataA(s_logisimBus227[10]),
.dataB(s_logisimBus283[10]),
.result(s_logisimNet366));
FullAdder
#(.extendedBits(2))
ARITH_2
(.carryIn(s_logisimBus443[11]),
.carryOut(s_logisimNet35),
.dataA(s_logisimBus227[11]),
.dataB(s_logisimBus283[11]),
.result(s_logisimNet296));
FullAdder
#(.extendedBits(2))
ARITH_3
(.carryIn(s_logisimBus443[12]),
.carryOut(s_logisimNet245),
.dataA(s_logisimBus227[12]),
.dataB(s_logisimBus283[12]),
.result(s_logisimNet213));
FullAdder
#(.extendedBits(2))
ARITH_4
(.carryIn(s_logisimBus443[13]),
.carryOut(s_logisimNet159),
.dataA(s_logisimBus227[13]),
.dataB(s_logisimBus283[13]),
.result(s_logisimNet124));
FullAdder
#(.extendedBits(2))
ARITH_5
(.carryIn(s_logisimBus443[14]),
.carryOut(s_logisimNet62),
.dataA(s_logisimBus227[14]),
.dataB(s_logisimBus283[14]),
.result(s_logisimNet14));
FullAdder
#(.extendedBits(2))
ARITH_6
(.carryIn(s_logisimBus443[15]),
.carryOut(s_logisimNet110),
.dataA(s_logisimBus227[15]),
.dataB(s_logisimBus283[15]),
.result(s_logisimNet390));
FullAdder
#(.extendedBits(2))
ARITH_7
(.carryIn(s_logisimBus443[16]),
.carryOut(s_logisimNet75),
.dataA(s_logisimBus227[16]),
.dataB(s_logisimBus283[16]),
.result(s_logisimNet320));
FullAdder
#(.extendedBits(2))
ARITH_8
(.carryIn(s_logisimBus443[17]),
.carryOut(s_logisimNet276),
.dataA(s_logisimBus227[17]),
.dataB(s_logisimBus283[17]),
.result(s_logisimNet243));
FullAdder
#(.extendedBits(2))
ARITH_9
(.carryIn(s_logisimBus443[18]),
.carryOut(s_logisimNet191),
.dataA(s_logisimBus227[18]),
.dataB(s_logisimBus283[18]),
.result(s_logisimNet158));
FullAdder
#(.extendedBits(2))
ARITH_10
(.carryIn(s_logisimBus443[19]),
.carryOut(s_logisimNet98),
.dataA(s_logisimBus227[19]),
.dataB(s_logisimBus283[19]),
.result(s_logisimNet57));
FullAdder
#(.extendedBits(2))
ARITH_11
(.carryIn(s_logisimBus443[20]),
.carryOut(s_logisimNet139),
.dataA(s_logisimBus227[20]),
.dataB(s_logisimBus283[20]),
.result(s_logisimNet412));
FullAdder
#(.extendedBits(2))
ARITH_12
(.carryIn(s_logisimBus443[21]),
.carryOut(s_logisimNet37),
.dataA(s_logisimBus227[21]),
.dataB(s_logisimBus283[21]),
.result(s_logisimNet345));
FullAdder
#(.extendedBits(2))
ARITH_13
(.carryIn(s_logisimBus443[22]),
.carryOut(s_logisimNet9),
.dataA(s_logisimBus227[22]),
.dataB(s_logisimBus283[22]),
.result(s_logisimNet270));
FullAdder
#(.extendedBits(2))
ARITH_14
(.carryIn(s_logisimBus443[23]),
.carryOut(s_logisimNet219),
.dataA(s_logisimBus227[23]),
.dataB(s_logisimBus283[23]),
.result(s_logisimNet184));
FullAdder
#(.extendedBits(2))
ARITH_15
(.carryIn(s_logisimBus443[24]),
.carryOut(s_logisimNet130),
.dataA(s_logisimBus227[24]),
.dataB(s_logisimBus283[24]),
.result(s_logisimNet92));
FullAdder
#(.extendedBits(2))
ARITH_16
(.carryIn(s_logisimBus443[25]),
.carryOut(s_logisimNet20),
.dataA(s_logisimBus227[25]),
.dataB(s_logisimBus283[25]),
.result(s_logisimNet430));
FullAdder
#(.extendedBits(2))
ARITH_17
(.carryIn(s_logisimBus443[26]),
.carryOut(s_logisimNet76),
.dataA(s_logisimBus227[26]),
.dataB(s_logisimBus283[26]),
.result(s_logisimNet367));
FullAdder
#(.extendedBits(2))
ARITH_18
(.carryIn(s_logisimBus443[1]),
.carryOut(s_logisimNet272),
.dataA(s_logisimBus227[1]),
.dataB(s_logisimBus283[1]),
.result(s_logisimNet241));
FullAdder
#(.extendedBits(2))
ARITH_19
(.carryIn(s_logisimBus443[27]),
.carryOut(s_logisimNet28),
.dataA(s_logisimBus227[27]),
.dataB(s_logisimBus283[27]),
.result(s_logisimNet297));
FullAdder
#(.extendedBits(2))
ARITH_20
(.carryIn(s_logisimBus443[28]),
.carryOut(s_logisimNet249),
.dataA(s_logisimBus227[28]),
.dataB(s_logisimBus283[28]),
.result(s_logisimNet214));
FullAdder
#(.extendedBits(2))
ARITH_21
(.carryIn(s_logisimBus443[29]),
.carryOut(s_logisimNet164),
.dataA(s_logisimBus227[29]),
.dataB(s_logisimBus283[29]),
.result(s_logisimNet125));
FullAdder
#(.extendedBits(2))
ARITH_22
(.carryIn(s_logisimBus443[30]),
.carryOut(s_logisimNet63),
.dataA(s_logisimBus227[30]),
.dataB(s_logisimBus283[30]),
.result(s_logisimNet17));
FullAdder
#(.extendedBits(2))
ARITH_23
(.carryIn(s_logisimBus443[31]),
.carryOut(s_logisimNet108),
.dataA(s_logisimBus227[31]),
.dataB(s_logisimBus283[31]),
.result(s_logisimNet393));
FullAdder
#(.extendedBits(2))
ARITH_24
(.carryIn(s_logisimBus443[32]),
.carryOut(s_logisimNet69),
.dataA(s_logisimBus227[32]),
.dataB(s_logisimBus283[32]),
.result(s_logisimNet323));
FullAdder
#(.extendedBits(2))
ARITH_25
(.carryIn(s_logisimBus443[33]),
.carryOut(s_logisimNet277),
.dataA(s_logisimBus227[33]),
.dataB(s_logisimBus283[33]),
.result(s_logisimNet246));
FullAdder
#(.extendedBits(2))
ARITH_26
(.carryIn(s_logisimBus443[34]),
.carryOut(s_logisimNet192),
.dataA(s_logisimBus227[34]),
.dataB(s_logisimBus283[34]),
.result(s_logisimNet160));
FullAdder
#(.extendedBits(2))
ARITH_27
(.carryIn(s_logisimBus443[35]),
.carryOut(s_logisimNet99),
.dataA(s_logisimBus227[35]),
.dataB(s_logisimBus283[35]),
.result(s_logisimNet58));
FullAdder
#(.extendedBits(2))
ARITH_28
(.carryIn(s_logisimBus443[36]),
.carryOut(s_logisimNet140),
.dataA(s_logisimBus227[36]),
.dataB(s_logisimBus283[36]),
.result(s_logisimNet414));
FullAdder
#(.extendedBits(2))
ARITH_29
(.carryIn(s_logisimBus443[2]),
.carryOut(s_logisimNet187),
.dataA(s_logisimBus227[2]),
.dataB(s_logisimBus283[2]),
.result(s_logisimNet156));
FullAdder
#(.extendedBits(2))
ARITH_30
(.carryIn(s_logisimBus443[37]),
.carryOut(s_logisimNet38),
.dataA(s_logisimBus227[37]),
.dataB(s_logisimBus283[37]),
.result(s_logisimNet347));
FullAdder
#(.extendedBits(2))
ARITH_31
(.carryIn(s_logisimBus443[38]),
.carryOut(s_logisimNet6),
.dataA(s_logisimBus227[38]),
.dataB(s_logisimBus283[38]),
.result(s_logisimNet273));
FullAdder
#(.extendedBits(2))
ARITH_32
(.carryIn(s_logisimBus443[39]),
.carryOut(s_logisimNet211),
.dataA(s_logisimBus227[39]),
.dataB(s_logisimBus283[39]),
.result(s_logisimNet188));
FullAdder
#(.extendedBits(2))
ARITH_33
(.carryIn(s_logisimBus443[40]),
.carryOut(s_logisimNet122),
.dataA(s_logisimBus227[40]),
.dataB(s_logisimBus283[40]),
.result(s_logisimNet96));
FullAdder
#(.extendedBits(2))
ARITH_34
(.carryIn(s_logisimBus443[41]),
.carryOut(s_logisimNet12),
.dataA(s_logisimBus227[41]),
.dataB(s_logisimBus283[41]),
.result(s_logisimNet433));
FullAdder
#(.extendedBits(2))
ARITH_35
(.carryIn(s_logisimBus443[42]),
.carryOut(s_logisimNet77),
.dataA(s_logisimBus227[42]),
.dataB(s_logisimBus283[42]),
.result(s_logisimNet369));
FullAdder
#(.extendedBits(2))
ARITH_36
(.carryIn(s_logisimBus443[43]),
.carryOut(s_logisimNet29),
.dataA(s_logisimBus227[43]),
.dataB(s_logisimBus283[43]),
.result(s_logisimNet299));
FullAdder
#(.extendedBits(2))
ARITH_37
(.carryIn(s_logisimBus443[44]),
.carryOut(s_logisimNet240),
.dataA(s_logisimBus227[44]),
.dataB(s_logisimBus283[44]),
.result(s_logisimNet217));
FullAdder
#(.extendedBits(2))
ARITH_38
(.carryIn(s_logisimBus443[45]),
.carryOut(s_logisimNet155),
.dataA(s_logisimBus227[45]),
.dataB(s_logisimBus283[45]),
.result(s_logisimNet128));
FullAdder
#(.extendedBits(2))
ARITH_39
(.carryIn(s_logisimBus443[46]),
.carryOut(s_logisimNet54),
.dataA(s_logisimBus227[46]),
.dataB(s_logisimBus283[46]),
.result(s_logisimNet18));
FullAdder
#(.extendedBits(2))
ARITH_40
(.carryIn(s_logisimBus443[3]),
.carryOut(s_logisimNet95),
.dataA(s_logisimBus227[3]),
.dataB(s_logisimBus283[3]),
.result(s_logisimNet55));
FullAdder
#(.extendedBits(2))
ARITH_41
(.carryIn(s_logisimBus443[47]),
.carryOut(s_logisimNet109),
.dataA(s_logisimBus227[47]),
.dataB(s_logisimBus283[47]),
.result(s_logisimNet394));
FullAdder
#(.extendedBits(2))
ARITH_42
(.carryIn(s_logisimBus443[48]),
.carryOut(s_logisimNet70),
.dataA(s_logisimBus227[48]),
.dataB(s_logisimBus283[48]),
.result(s_logisimNet324));
FullAdder
#(.extendedBits(2))
ARITH_43
(.carryIn(s_logisimBus443[49]),
.carryOut(s_logisimNet268),
.dataA(s_logisimBus227[49]),
.dataB(s_logisimBus283[49]),
.result(s_logisimNet247));
FullAdder
#(.extendedBits(2))
ARITH_44
(.carryIn(s_logisimBus443[50]),
.carryOut(s_logisimNet183),
.dataA(s_logisimBus227[50]),
.dataB(s_logisimBus283[50]),
.result(s_logisimNet161));
FullAdder
#(.extendedBits(2))
ARITH_45
(.carryIn(s_logisimBus443[51]),
.carryOut(s_logisimNet91),
.dataA(s_logisimBus227[51]),
.dataB(s_logisimBus283[51]),
.result(s_logisimNet59));
FullAdder
#(.extendedBits(2))
ARITH_46
(.carryIn(s_logisimBus443[52]),
.carryOut(s_logisimNet141),
.dataA(s_logisimBus227[52]),
.dataB(s_logisimBus283[52]),
.result(s_logisimNet415));
FullAdder
#(.extendedBits(2))
ARITH_47
(.carryIn(s_logisimBus443[53]),
.carryOut(s_logisimNet39),
.dataA(s_logisimBus227[53]),
.dataB(s_logisimBus283[53]),
.result(s_logisimNet350));
FullAdder
#(.extendedBits(2))
ARITH_48
(.carryIn(s_logisimBus443[54]),
.carryOut(s_logisimNet7),
.dataA(s_logisimBus227[54]),
.dataB(s_logisimBus283[54]),
.result(s_logisimNet278));
FullAdder
#(.extendedBits(2))
ARITH_49
(.carryIn(s_logisimBus443[55]),
.carryOut(s_logisimNet212),
.dataA(s_logisimBus227[55]),
.dataB(s_logisimBus283[55]),
.result(s_logisimNet193));
FullAdder
#(.extendedBits(2))
ARITH_50
(.carryIn(s_logisimBus443[56]),
.carryOut(s_logisimNet123),
.dataA(s_logisimBus227[56]),
.dataB(s_logisimBus283[56]),
.result(s_logisimNet100));
FullAdder
#(.extendedBits(2))
ARITH_51
(.carryIn(s_logisimBus443[4]),
.carryOut(s_logisimNet143),
.dataA(s_logisimBus227[4]),
.dataB(s_logisimBus283[4]),
.result(s_logisimNet411));
FullAdder
#(.extendedBits(2))
ARITH_52
(.carryIn(s_logisimBus443[57]),
.carryOut(s_logisimNet13),
.dataA(s_logisimBus227[57]),
.dataB(s_logisimBus283[57]),
.result(s_logisimNet435));
FullAdder
#(.extendedBits(2))
ARITH_53
(.carryIn(s_logisimBus443[58]),
.carryOut(s_logisimNet78),
.dataA(s_logisimBus227[58]),
.dataB(s_logisimBus283[58]),
.result(s_logisimNet371));
FullAdder
#(.extendedBits(2))
ARITH_54
(.carryIn(s_logisimBus443[59]),
.carryOut(s_logisimNet30),
.dataA(s_logisimBus227[59]),
.dataB(s_logisimBus283[59]),
.result(s_logisimNet301));
FullAdder
#(.extendedBits(2))
ARITH_55
(.carryIn(s_logisimBus443[60]),
.carryOut(s_logisimNet242),
.dataA(s_logisimBus227[60]),
.dataB(s_logisimBus283[60]),
.result(s_logisimNet220));
FullAdder
#(.extendedBits(2))
ARITH_56
(.carryIn(s_logisimBus443[61]),
.carryOut(s_logisimNet157),
.dataA(s_logisimBus227[61]),
.dataB(s_logisimBus283[61]),
.result(s_logisimNet131));
FullAdder
#(.extendedBits(2))
ARITH_57
(.carryIn(s_logisimBus443[62]),
.carryOut(s_logisimNet56),
.dataA(s_logisimBus227[62]),
.dataB(s_logisimBus283[62]),
.result(s_logisimNet21));
FullAdder
#(.extendedBits(2))
ARITH_58
(.carryIn(s_logisimBus443[63]),
.carryOut(),
.dataA(s_logisimBus227[63]),
.dataB(s_logisimBus283[63]),
.result(s_logisimNet396));
FullAdder
#(.extendedBits(2))
ARITH_59
(.carryIn(s_logisimBus443[5]),
.carryOut(s_logisimNet41),
.dataA(s_logisimBus227[5]),
.dataB(s_logisimBus283[5]),
.result(s_logisimNet344));
FullAdder
#(.extendedBits(2))
ARITH_60
(.carryIn(s_logisimBus443[6]),
.carryOut(s_logisimNet8),
.dataA(s_logisimBus227[6]),
.dataB(s_logisimBus283[6]),
.result(s_logisimNet269));
FullAdder
#(.extendedBits(2))
ARITH_61
(.carryIn(s_logisimBus443[7]),
.carryOut(s_logisimNet216),
.dataA(s_logisimBus227[7]),
.dataB(s_logisimBus283[7]),
.result(s_logisimNet185));
FullAdder
#(.extendedBits(2))
ARITH_62
(.carryIn(s_logisimBus443[8]),
.carryOut(s_logisimNet127),
.dataA(s_logisimBus227[8]),
.dataB(s_logisimBus283[8]),
.result(s_logisimNet93));
FullAdder
#(.extendedBits(2))
ARITH_63
(.carryIn(s_logisimBus443[9]),
.carryOut(s_logisimNet15),
.dataA(s_logisimBus227[9]),
.dataB(s_logisimBus283[9]),
.result(s_logisimNet431));
FullAdder
#(.extendedBits(2))
ARITH_64
(.carryIn(s_logisimNet138),
.carryOut(s_logisimNet42),
.dataA(s_logisimNet15),
.dataB(s_logisimNet366),
.result(s_logisimBus448[10]));
FullAdder
#(.extendedBits(2))
ARITH_65
(.carryIn(s_logisimNet42),
.carryOut(s_logisimNet403),
.dataA(s_logisimNet79),
.dataB(s_logisimNet296),
.result(s_logisimBus448[11]));
FullAdder
#(.extendedBits(2))
ARITH_66
(.carryIn(s_logisimNet403),
.carryOut(s_logisimNet332),
.dataA(s_logisimNet35),
.dataB(s_logisimNet213),
.result(s_logisimBus448[12]));
FullAdder
#(.extendedBits(2))
ARITH_67
(.carryIn(s_logisimNet332),
.carryOut(s_logisimNet256),
.dataA(s_logisimNet245),
.dataB(s_logisimNet124),
.result(s_logisimBus448[13]));
FullAdder
#(.extendedBits(2))
ARITH_68
(.carryIn(s_logisimNet256),
.carryOut(s_logisimNet171),
.dataA(s_logisimNet159),
.dataB(s_logisimNet14),
.result(s_logisimBus448[14]));
FullAdder
#(.extendedBits(2))
ARITH_69
(.carryIn(s_logisimNet171),
.carryOut(s_logisimNet80),
.dataA(s_logisimNet62),
.dataB(s_logisimNet390),
.result(s_logisimBus448[15]));
FullAdder
#(.extendedBits(2))
ARITH_70
(.carryIn(s_logisimBus443[0]),
.carryOut(s_logisimNet422),
.dataA(s_logisimBus227[0]),
.dataB(s_logisimBus283[0]),
.result(s_logisimBus448[0]));
FullAdder
#(.extendedBits(2))
ARITH_71
(.carryIn(s_logisimNet80),
.carryOut(s_logisimNet423),
.dataA(s_logisimNet110),
.dataB(s_logisimNet320),
.result(s_logisimBus448[16]));
FullAdder
#(.extendedBits(2))
ARITH_72
(.carryIn(s_logisimNet423),
.carryOut(s_logisimNet356),
.dataA(s_logisimNet75),
.dataB(s_logisimNet243),
.result(s_logisimBus448[17]));
FullAdder
#(.extendedBits(2))
ARITH_73
(.carryIn(s_logisimNet356),
.carryOut(s_logisimNet285),
.dataA(s_logisimNet276),
.dataB(s_logisimNet158),
.result(s_logisimBus448[18]));
FullAdder
#(.extendedBits(2))
ARITH_74
(.carryIn(s_logisimNet285),
.carryOut(s_logisimNet200),
.dataA(s_logisimNet191),
.dataB(s_logisimNet57),
.result(s_logisimBus448[19]));
FullAdder
#(.extendedBits(2))
ARITH_75
(.carryIn(s_logisimNet200),
.carryOut(s_logisimNet111),
.dataA(s_logisimNet98),
.dataB(s_logisimNet412),
.result(s_logisimBus448[20]));
FullAdder
#(.extendedBits(2))
ARITH_76
(.carryIn(s_logisimNet111),
.carryOut(s_logisimNet445),
.dataA(s_logisimNet139),
.dataB(s_logisimNet345),
.result(s_logisimBus448[21]));
FullAdder
#(.extendedBits(2))
ARITH_77
(.carryIn(s_logisimNet445),
.carryOut(s_logisimNet379),
.dataA(s_logisimNet37),
.dataB(s_logisimNet270),
.result(s_logisimBus448[22]));
FullAdder
#(.extendedBits(2))
ARITH_78
(.carryIn(s_logisimNet379),
.carryOut(s_logisimNet310),
.dataA(s_logisimNet9),
.dataB(s_logisimNet184),
.result(s_logisimBus448[23]));
FullAdder
#(.extendedBits(2))
ARITH_79
(.carryIn(s_logisimNet310),
.carryOut(s_logisimNet230),
.dataA(s_logisimNet219),
.dataB(s_logisimNet92),
.result(s_logisimBus448[24]));
FullAdder
#(.extendedBits(2))
ARITH_80
(.carryIn(s_logisimNet230),
.carryOut(s_logisimNet144),
.dataA(s_logisimNet130),
.dataB(s_logisimNet430),
.result(s_logisimBus448[25]));
FullAdder
#(.extendedBits(2))
ARITH_81
(.carryIn(s_logisimNet422),
.carryOut(s_logisimNet355),
.dataA(s_logisimNet444),
.dataB(s_logisimNet241),
.result(s_logisimBus448[1]));
FullAdder
#(.extendedBits(2))
ARITH_82
(.carryIn(s_logisimNet144),
.carryOut(s_logisimNet43),
.dataA(s_logisimNet20),
.dataB(s_logisimNet367),
.result(s_logisimBus448[26]));
FullAdder
#(.extendedBits(2))
ARITH_83
(.carryIn(s_logisimNet43),
.carryOut(s_logisimNet404),
.dataA(s_logisimNet76),
.dataB(s_logisimNet297),
.result(s_logisimBus448[27]));
FullAdder
#(.extendedBits(2))
ARITH_84
(.carryIn(s_logisimNet404),
.carryOut(s_logisimNet333),
.dataA(s_logisimNet28),
.dataB(s_logisimNet214),
.result(s_logisimBus448[28]));
FullAdder
#(.extendedBits(2))
ARITH_85
(.carryIn(s_logisimNet333),
.carryOut(s_logisimNet257),
.dataA(s_logisimNet249),
.dataB(s_logisimNet125),
.result(s_logisimBus448[29]));
FullAdder
#(.extendedBits(2))
ARITH_86
(.carryIn(s_logisimNet257),
.carryOut(s_logisimNet172),
.dataA(s_logisimNet164),
.dataB(s_logisimNet17),
.result(s_logisimBus448[30]));
FullAdder
#(.extendedBits(2))
ARITH_87
(.carryIn(s_logisimNet172),
.carryOut(s_logisimNet81),
.dataA(s_logisimNet63),
.dataB(s_logisimNet393),
.result(s_logisimBus448[31]));
FullAdder
#(.extendedBits(2))
ARITH_88
(.carryIn(s_logisimNet81),
.carryOut(s_logisimNet424),
.dataA(s_logisimNet108),
.dataB(s_logisimNet323),
.result(s_logisimBus448[32]));
FullAdder
#(.extendedBits(2))
ARITH_89
(.carryIn(s_logisimNet424),
.carryOut(s_logisimNet357),
.dataA(s_logisimNet69),
.dataB(s_logisimNet246),
.result(s_logisimBus448[33]));
FullAdder
#(.extendedBits(2))
ARITH_90
(.carryIn(s_logisimNet357),
.carryOut(s_logisimNet286),
.dataA(s_logisimNet277),
.dataB(s_logisimNet160),
.result(s_logisimBus448[34]));
FullAdder
#(.extendedBits(2))
ARITH_91
(.carryIn(s_logisimNet286),
.carryOut(s_logisimNet201),
.dataA(s_logisimNet192),
.dataB(s_logisimNet58),
.result(s_logisimBus448[35]));
FullAdder
#(.extendedBits(2))
ARITH_92
(.carryIn(s_logisimNet355),
.carryOut(s_logisimNet284),
.dataA(s_logisimNet272),
.dataB(s_logisimNet156),
.result(s_logisimBus448[2]));
FullAdder
#(.extendedBits(2))
ARITH_93
(.carryIn(s_logisimNet201),
.carryOut(s_logisimNet112),
.dataA(s_logisimNet99),
.dataB(s_logisimNet414),
.result(s_logisimBus448[36]));
FullAdder
#(.extendedBits(2))
ARITH_94
(.carryIn(s_logisimNet112),
.carryOut(s_logisimNet446),
.dataA(s_logisimNet140),
.dataB(s_logisimNet347),
.result(s_logisimBus448[37]));
FullAdder
#(.extendedBits(2))
ARITH_95
(.carryIn(s_logisimNet446),
.carryOut(s_logisimNet380),
.dataA(s_logisimNet38),
.dataB(s_logisimNet273),
.result(s_logisimBus448[38]));
FullAdder
#(.extendedBits(2))
ARITH_96
(.carryIn(s_logisimNet380),
.carryOut(s_logisimNet311),
.dataA(s_logisimNet6),
.dataB(s_logisimNet188),
.result(s_logisimBus448[39]));
FullAdder
#(.extendedBits(2))
ARITH_97
(.carryIn(s_logisimNet311),
.carryOut(s_logisimNet231),
.dataA(s_logisimNet211),
.dataB(s_logisimNet96),
.result(s_logisimBus448[40]));
FullAdder
#(.extendedBits(2))
ARITH_98
(.carryIn(s_logisimNet231),
.carryOut(s_logisimNet145),
.dataA(s_logisimNet122),
.dataB(s_logisimNet433),
.result(s_logisimBus448[41]));
FullAdder
#(.extendedBits(2))
ARITH_99
(.carryIn(s_logisimNet145),
.carryOut(s_logisimNet44),
.dataA(s_logisimNet12),
.dataB(s_logisimNet369),
.result(s_logisimBus448[42]));
FullAdder
#(.extendedBits(2))
ARITH_100
(.carryIn(s_logisimNet44),
.carryOut(s_logisimNet405),
.dataA(s_logisimNet77),
.dataB(s_logisimNet299),
.result(s_logisimBus448[43]));
FullAdder
#(.extendedBits(2))
ARITH_101
(.carryIn(s_logisimNet405),
.carryOut(s_logisimNet334),
.dataA(s_logisimNet29),
.dataB(s_logisimNet217),
.result(s_logisimBus448[44]));
FullAdder
#(.extendedBits(2))
ARITH_102
(.carryIn(s_logisimNet334),
.carryOut(s_logisimNet258),
.dataA(s_logisimNet240),
.dataB(s_logisimNet128),
.result(s_logisimBus448[45]));
FullAdder
#(.extendedBits(2))
ARITH_103
(.carryIn(s_logisimNet284),
.carryOut(s_logisimNet199),
.dataA(s_logisimNet187),
.dataB(s_logisimNet55),
.result(s_logisimBus448[3]));
FullAdder
#(.extendedBits(2))
ARITH_104
(.carryIn(s_logisimNet258),
.carryOut(s_logisimNet173),
.dataA(s_logisimNet155),
.dataB(s_logisimNet18),
.result(s_logisimBus448[46]));
FullAdder
#(.extendedBits(2))
ARITH_105
(.carryIn(s_logisimNet173),
.carryOut(s_logisimNet82),
.dataA(s_logisimNet54),
.dataB(s_logisimNet394),
.result(s_logisimBus448[47]));
FullAdder
#(.extendedBits(2))
ARITH_106
(.carryIn(s_logisimNet82),
.carryOut(s_logisimNet425),
.dataA(s_logisimNet109),
.dataB(s_logisimNet324),
.result(s_logisimBus448[48]));
FullAdder
#(.extendedBits(2))
ARITH_107
(.carryIn(s_logisimNet425),
.carryOut(s_logisimNet358),
.dataA(s_logisimNet70),
.dataB(s_logisimNet247),
.result(s_logisimBus448[49]));
FullAdder
#(.extendedBits(2))
ARITH_108
(.carryIn(s_logisimNet358),
.carryOut(s_logisimNet287),
.dataA(s_logisimNet268),
.dataB(s_logisimNet161),
.result(s_logisimBus448[50]));
FullAdder
#(.extendedBits(2))
ARITH_109
(.carryIn(s_logisimNet287),
.carryOut(s_logisimNet202),
.dataA(s_logisimNet183),
.dataB(s_logisimNet59),
.result(s_logisimBus448[51]));
FullAdder
#(.extendedBits(2))
ARITH_110
(.carryIn(s_logisimNet202),
.carryOut(s_logisimNet113),
.dataA(s_logisimNet91),
.dataB(s_logisimNet415),
.result(s_logisimBus448[52]));
FullAdder
#(.extendedBits(2))
ARITH_111
(.carryIn(s_logisimNet113),
.carryOut(s_logisimNet447),
.dataA(s_logisimNet141),
.dataB(s_logisimNet350),
.result(s_logisimBus448[53]));
FullAdder
#(.extendedBits(2))
ARITH_112
(.carryIn(s_logisimNet447),
.carryOut(s_logisimNet381),
.dataA(s_logisimNet39),
.dataB(s_logisimNet278),
.result(s_logisimBus448[54]));
FullAdder
#(.extendedBits(2))
ARITH_113
(.carryIn(s_logisimNet381),
.carryOut(s_logisimNet309),
.dataA(s_logisimNet7),
.dataB(s_logisimNet193),
.result(s_logisimBus448[55]));
FullAdder
#(.extendedBits(2))
ARITH_114
(.carryIn(s_logisimNet199),
.carryOut(s_logisimNet107),
.dataA(s_logisimNet95),
.dataB(s_logisimNet411),
.result(s_logisimBus448[4]));
FullAdder
#(.extendedBits(2))
ARITH_115
(.carryIn(s_logisimNet309),
.carryOut(s_logisimNet229),
.dataA(s_logisimNet212),
.dataB(s_logisimNet100),
.result(s_logisimBus448[56]));
FullAdder
#(.extendedBits(2))
ARITH_116
(.carryIn(s_logisimNet229),
.carryOut(s_logisimNet142),
.dataA(s_logisimNet123),
.dataB(s_logisimNet435),
.result(s_logisimBus448[57]));
FullAdder
#(.extendedBits(2))
ARITH_117
(.carryIn(s_logisimNet142),
.carryOut(s_logisimNet40),
.dataA(s_logisimNet13),
.dataB(s_logisimNet371),
.result(s_logisimBus448[58]));
FullAdder
#(.extendedBits(2))
ARITH_118
(.carryIn(s_logisimNet40),
.carryOut(s_logisimNet402),
.dataA(s_logisimNet78),
.dataB(s_logisimNet301),
.result(s_logisimBus448[59]));
FullAdder
#(.extendedBits(2))
ARITH_119
(.carryIn(s_logisimNet402),
.carryOut(s_logisimNet331),
.dataA(s_logisimNet30),
.dataB(s_logisimNet220),
.result(s_logisimBus448[60]));
FullAdder
#(.extendedBits(2))
ARITH_120
(.carryIn(s_logisimNet331),
.carryOut(s_logisimNet255),
.dataA(s_logisimNet242),
.dataB(s_logisimNet131),
.result(s_logisimBus448[61]));
FullAdder
#(.extendedBits(2))
ARITH_121
(.carryIn(s_logisimNet255),
.carryOut(s_logisimNet170),
.dataA(s_logisimNet157),
.dataB(s_logisimNet21),
.result(s_logisimBus448[62]));
FullAdder
#(.extendedBits(2))
ARITH_122
(.carryIn(s_logisimNet170),
.carryOut(),
.dataA(s_logisimNet56),
.dataB(s_logisimNet396),
.result(s_logisimBus448[63]));
FullAdder
#(.extendedBits(2))
ARITH_123
(.carryIn(s_logisimNet107),
.carryOut(s_logisimNet442),
.dataA(s_logisimNet143),
.dataB(s_logisimNet344),
.result(s_logisimBus448[5]));
FullAdder
#(.extendedBits(2))
ARITH_124
(.carryIn(s_logisimNet442),
.carryOut(s_logisimNet378),
.dataA(s_logisimNet41),
.dataB(s_logisimNet269),
.result(s_logisimBus448[6]));
FullAdder
#(.extendedBits(2))
ARITH_125
(.carryIn(s_logisimNet378),
.carryOut(s_logisimNet308),
.dataA(s_logisimNet8),
.dataB(s_logisimNet185),
.result(s_logisimBus448[7]));
FullAdder
#(.extendedBits(2))
ARITH_126
(.carryIn(s_logisimNet308),
.carryOut(s_logisimNet228),
.dataA(s_logisimNet216),
.dataB(s_logisimNet93),
.result(s_logisimBus448[8]));
FullAdder
#(.extendedBits(2))
ARITH_127
(.carryIn(s_logisimNet228),
.carryOut(s_logisimNet138),
.dataA(s_logisimNet127),
.dataB(s_logisimNet431),
.result(s_logisimBus448[9]));
endmodule