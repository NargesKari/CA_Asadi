/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
SLL1
**
**
**
*****************************************************************************/
module
SLL1(
a,
b,
output1
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[31:0]
b;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[63:0]
output1;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[63:0]
s_logisimBus0;
wire
[4:0]
s_logisimBus1;
wire
[5:0]
s_logisimBus10;
wire
[4:0]
s_logisimBus11;
wire
[63:0]
s_logisimBus12;
wire
[31:0]
s_logisimBus14;
wire
[5:0]
s_logisimBus16;
wire
[63:0]
s_logisimBus17;
wire
[63:0]
s_logisimBus18;
wire
[31:0]
s_logisimBus2;
wire
[63:0]
s_logisimBus3;
wire
[5:0]
s_logisimBus4;
wire
[4:0]
s_logisimBus5;
wire
[63:0]
s_logisimBus6;
wire
[31:0]
s_logisimBus7;
wire
s_logisimNet15;
wire
s_logisimNet19;
wire
s_logisimNet20;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
wiring
is
defined
**
*******************************************************************************/
assign
s_logisimBus10[0]
=
s_logisimBus5[0];
assign
s_logisimBus10[1]
=
s_logisimBus5[1];
assign
s_logisimBus10[2]
=
s_logisimBus5[2];
assign
s_logisimBus10[3]
=
s_logisimBus5[3];
assign
s_logisimBus10[4]
=
s_logisimBus5[4];
assign
s_logisimBus1[0]
=
s_logisimBus2[0];
assign
s_logisimBus1[1]
=
s_logisimBus2[1];
assign
s_logisimBus1[2]
=
s_logisimBus2[2];
assign
s_logisimBus1[3]
=
s_logisimBus2[3];
assign
s_logisimBus1[4]
=
s_logisimBus2[4];
assign
s_logisimBus4[0]
=
s_logisimBus1[0];
assign
s_logisimBus4[1]
=
s_logisimBus1[1];
assign
s_logisimBus4[2]
=
s_logisimBus1[2];
assign
s_logisimBus4[3]
=
s_logisimBus1[3];
assign
s_logisimBus4[4]
=
s_logisimBus1[4];
assign
s_logisimBus5[0]
=
s_logisimBus14[0];
assign
s_logisimBus5[1]
=
s_logisimBus14[1];
assign
s_logisimBus5[2]
=
s_logisimBus14[2];
assign
s_logisimBus5[3]
=
s_logisimBus14[3];
assign
s_logisimBus5[4]
=
s_logisimBus14[4];
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus2[31:0]
=
b;
assign
s_logisimBus6[31:0]
=
a;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
output1
=
s_logisimBus0[63:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus6[63:32]
=
32'h00000000;
assign
s_logisimBus16[5:0]
=
{2'b00,
4'h1};
assign
s_logisimBus7[31:0]
=
32'h00000001;
assign
s_logisimBus4[5]
=
1'b0;
assign
s_logisimBus10[5]
=
1'b0;
assign
s_logisimBus11[4:0]
=
{1'b0,
4'h0};
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_1
(.enable(1'b1),
.muxIn_0(s_logisimBus12[63:0]),
.muxIn_1(s_logisimBus18[63:0]),
.muxOut(s_logisimBus17[63:0]),
.sel(s_logisimBus2[0]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus17[63:0]),
.muxIn_1(s_logisimBus6[63:0]),
.muxOut(s_logisimBus0[63:0]),
.sel(s_logisimNet15));
Shifter_64_bit
#(.shifterMode(0))
ARITH_3
(.dataA(s_logisimBus6[63:0]),
.result(s_logisimBus3[63:0]),
.shiftAmount(s_logisimBus16[5:0]));
Subtractor
#(.extendedBits(33),
.nrOfBits(32))
ARITH_4
(.borrowIn(1'b0),
.borrowOut(),
.dataA(s_logisimBus2[31:0]),
.dataB(s_logisimBus7[31:0]),
.result(s_logisimBus14[31:0]));
Shifter_64_bit
#(.shifterMode(0))
ARITH_5
(.dataA(s_logisimBus6[63:0]),
.result(s_logisimBus18[63:0]),
.shiftAmount(s_logisimBus4[5:0]));
Shifter_64_bit
#(.shifterMode(0))
ARITH_6
(.dataA(s_logisimBus3[63:0]),
.result(s_logisimBus12[63:0]),
.shiftAmount(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(5),
.twosComplement(1))
ARITH_7
(.aEqualsB(s_logisimNet15),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus1[4:0]),
.dataB(s_logisimBus11[4:0]));
endmodule