/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
ALU_SRA
**
**
**
*****************************************************************************/
module
ALU_SRA(
a,
b,
output1
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[31:0]
b;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[63:0]
output1;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[63:0]
s_logisimBus10;
wire
[63:0]
s_logisimBus12;
wire
[31:0]
s_logisimBus13;
wire
[5:0]
s_logisimBus14;
wire
[31:0]
s_logisimBus17;
wire
[63:0]
s_logisimBus18;
wire
[31:0]
s_logisimBus19;
wire
[31:0]
s_logisimBus2;
wire
[63:0]
s_logisimBus20;
wire
[63:0]
s_logisimBus21;
wire
[31:0]
s_logisimBus22;
wire
[31:0]
s_logisimBus23;
wire
[31:0]
s_logisimBus24;
wire
[5:0]
s_logisimBus25;
wire
[63:0]
s_logisimBus3;
wire
[63:0]
s_logisimBus5;
wire
[7:0]
s_logisimBus7;
wire
[31:0]
s_logisimBus9;
wire
s_logisimNet11;
wire
s_logisimNet15;
wire
s_logisimNet4;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
wiring
is
defined
**
*******************************************************************************/
assign
s_logisimBus20[0]
=
s_logisimBus2[0];
assign
s_logisimBus20[10]
=
s_logisimBus2[10];
assign
s_logisimBus20[11]
=
s_logisimBus2[11];
assign
s_logisimBus20[12]
=
s_logisimBus2[12];
assign
s_logisimBus20[13]
=
s_logisimBus2[13];
assign
s_logisimBus20[14]
=
s_logisimBus2[14];
assign
s_logisimBus20[15]
=
s_logisimBus2[15];
assign
s_logisimBus20[16]
=
s_logisimBus2[16];
assign
s_logisimBus20[17]
=
s_logisimBus2[17];
assign
s_logisimBus20[18]
=
s_logisimBus2[18];
assign
s_logisimBus20[19]
=
s_logisimBus2[19];
assign
s_logisimBus20[1]
=
s_logisimBus2[1];
assign
s_logisimBus20[20]
=
s_logisimBus2[20];
assign
s_logisimBus20[21]
=
s_logisimBus2[21];
assign
s_logisimBus20[22]
=
s_logisimBus2[22];
assign
s_logisimBus20[23]
=
s_logisimBus2[23];
assign
s_logisimBus20[24]
=
s_logisimBus2[24];
assign
s_logisimBus20[25]
=
s_logisimBus2[25];
assign
s_logisimBus20[26]
=
s_logisimBus2[26];
assign
s_logisimBus20[27]
=
s_logisimBus2[27];
assign
s_logisimBus20[28]
=
s_logisimBus2[28];
assign
s_logisimBus20[29]
=
s_logisimBus2[29];
assign
s_logisimBus20[2]
=
s_logisimBus2[2];
assign
s_logisimBus20[30]
=
s_logisimBus2[30];
assign
s_logisimBus20[31]
=
s_logisimBus2[31];
assign
s_logisimBus20[3]
=
s_logisimBus2[3];
assign
s_logisimBus20[4]
=
s_logisimBus2[4];
assign
s_logisimBus20[5]
=
s_logisimBus2[5];
assign
s_logisimBus20[6]
=
s_logisimBus2[6];
assign
s_logisimBus20[7]
=
s_logisimBus2[7];
assign
s_logisimBus20[8]
=
s_logisimBus2[8];
assign
s_logisimBus20[9]
=
s_logisimBus2[9];
assign
s_logisimBus2[0]
=
s_logisimBus10[0];
assign
s_logisimBus2[10]
=
s_logisimBus10[10];
assign
s_logisimBus2[11]
=
s_logisimBus10[11];
assign
s_logisimBus2[12]
=
s_logisimBus10[12];
assign
s_logisimBus2[13]
=
s_logisimBus10[13];
assign
s_logisimBus2[14]
=
s_logisimBus10[14];
assign
s_logisimBus2[15]
=
s_logisimBus10[15];
assign
s_logisimBus2[16]
=
s_logisimBus10[16];
assign
s_logisimBus2[17]
=
s_logisimBus10[17];
assign
s_logisimBus2[18]
=
s_logisimBus10[18];
assign
s_logisimBus2[19]
=
s_logisimBus10[19];
assign
s_logisimBus2[1]
=
s_logisimBus10[1];
assign
s_logisimBus2[20]
=
s_logisimBus10[20];
assign
s_logisimBus2[21]
=
s_logisimBus10[21];
assign
s_logisimBus2[22]
=
s_logisimBus10[22];
assign
s_logisimBus2[23]
=
s_logisimBus10[23];
assign
s_logisimBus2[24]
=
s_logisimBus10[24];
assign
s_logisimBus2[25]
=
s_logisimBus10[25];
assign
s_logisimBus2[26]
=
s_logisimBus10[26];
assign
s_logisimBus2[27]
=
s_logisimBus10[27];
assign
s_logisimBus2[28]
=
s_logisimBus10[28];
assign
s_logisimBus2[29]
=
s_logisimBus10[29];
assign
s_logisimBus2[2]
=
s_logisimBus10[2];
assign
s_logisimBus2[30]
=
s_logisimBus10[30];
assign
s_logisimBus2[31]
=
s_logisimBus10[31];
assign
s_logisimBus2[3]
=
s_logisimBus10[3];
assign
s_logisimBus2[4]
=
s_logisimBus10[4];
assign
s_logisimBus2[5]
=
s_logisimBus10[5];
assign
s_logisimBus2[6]
=
s_logisimBus10[6];
assign
s_logisimBus2[7]
=
s_logisimBus10[7];
assign
s_logisimBus2[8]
=
s_logisimBus10[8];
assign
s_logisimBus2[9]
=
s_logisimBus10[9];
assign
s_logisimBus9[16]
=
s_logisimBus7[0];
assign
s_logisimBus9[17]
=
s_logisimBus7[1];
assign
s_logisimBus9[18]
=
s_logisimBus7[2];
assign
s_logisimBus9[19]
=
s_logisimBus7[3];
assign
s_logisimBus9[20]
=
s_logisimBus7[4];
assign
s_logisimBus9[21]
=
s_logisimBus7[5];
assign
s_logisimBus9[22]
=
s_logisimBus7[6];
assign
s_logisimBus9[23]
=
s_logisimBus7[7];
assign
s_logisimBus9[24]
=
s_logisimBus7[0];
assign
s_logisimBus9[25]
=
s_logisimBus7[1];
assign
s_logisimBus9[26]
=
s_logisimBus7[2];
assign
s_logisimBus9[27]
=
s_logisimBus7[3];
assign
s_logisimBus9[28]
=
s_logisimBus7[4];
assign
s_logisimBus9[29]
=
s_logisimBus7[5];
assign
s_logisimBus9[30]
=
s_logisimBus7[6];
assign
s_logisimBus9[31]
=
s_logisimBus7[7];
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus17[31:0]
=
a;
assign
s_logisimBus19[31:0]
=
b;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
output1
=
s_logisimBus20[63:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus9[15:5]
=
{3'b000,
8'h00};
assign
s_logisimBus7[7:0]
=
8'h00;
assign
s_logisimBus9[0]
=
s_logisimBus19[0];
assign
s_logisimBus9[1]
=
s_logisimBus19[1];
assign
s_logisimBus9[2]
=
s_logisimBus19[2];
assign
s_logisimBus9[3]
=
s_logisimBus19[3];
assign
s_logisimBus9[4]
=
s_logisimBus19[4];
assign
s_logisimBus5[0]
=
s_logisimBus17[0];
assign
s_logisimBus5[1]
=
s_logisimBus17[1];
assign
s_logisimBus5[2]
=
s_logisimBus17[2];
assign
s_logisimBus5[3]
=
s_logisimBus17[3];
assign
s_logisimBus5[4]
=
s_logisimBus17[4];
assign
s_logisimBus5[5]
=
s_logisimBus17[5];
assign
s_logisimBus5[6]
=
s_logisimBus17[6];
assign
s_logisimBus5[7]
=
s_logisimBus17[7];
assign
s_logisimBus5[8]
=
s_logisimBus17[8];
assign
s_logisimBus5[9]
=
s_logisimBus17[9];
assign
s_logisimBus5[10]
=
s_logisimBus17[10];
assign
s_logisimBus5[11]
=
s_logisimBus17[11];
assign
s_logisimBus5[12]
=
s_logisimBus17[12];
assign
s_logisimBus5[13]
=
s_logisimBus17[13];
assign
s_logisimBus5[14]
=
s_logisimBus17[14];
assign
s_logisimBus5[15]
=
s_logisimBus17[15];
assign
s_logisimBus5[16]
=
s_logisimBus17[16];
assign
s_logisimBus5[17]
=
s_logisimBus17[17];
assign
s_logisimBus5[18]
=
s_logisimBus17[18];
assign
s_logisimBus5[19]
=
s_logisimBus17[19];
assign
s_logisimBus5[20]
=
s_logisimBus17[20];
assign
s_logisimBus5[21]
=
s_logisimBus17[21];
assign
s_logisimBus5[22]
=
s_logisimBus17[22];
assign
s_logisimBus5[23]
=
s_logisimBus17[23];
assign
s_logisimBus5[24]
=
s_logisimBus17[24];
assign
s_logisimBus5[25]
=
s_logisimBus17[25];
assign
s_logisimBus5[26]
=
s_logisimBus17[26];
assign
s_logisimBus5[27]
=
s_logisimBus17[27];
assign
s_logisimBus5[28]
=
s_logisimBus17[28];
assign
s_logisimBus5[29]
=
s_logisimBus17[29];
assign
s_logisimBus5[30]
=
s_logisimBus17[30];
assign
s_logisimBus5[31]
=
s_logisimBus17[31];
assign
s_logisimBus5[32]
=
s_logisimBus17[31];
assign
s_logisimBus5[33]
=
s_logisimBus17[31];
assign
s_logisimBus5[34]
=
s_logisimBus17[31];
assign
s_logisimBus5[35]
=
s_logisimBus17[31];
assign
s_logisimBus5[36]
=
s_logisimBus17[31];
assign
s_logisimBus5[37]
=
s_logisimBus17[31];
assign
s_logisimBus5[38]
=
s_logisimBus17[31];
assign
s_logisimBus5[39]
=
s_logisimBus17[31];
assign
s_logisimBus5[40]
=
s_logisimBus17[31];
assign
s_logisimBus5[41]
=
s_logisimBus17[31];
assign
s_logisimBus5[42]
=
s_logisimBus17[31];
assign
s_logisimBus5[43]
=
s_logisimBus17[31];
assign
s_logisimBus5[44]
=
s_logisimBus17[31];
assign
s_logisimBus5[45]
=
s_logisimBus17[31];
assign
s_logisimBus5[46]
=
s_logisimBus17[31];
assign
s_logisimBus5[47]
=
s_logisimBus17[31];
assign
s_logisimBus5[48]
=
s_logisimBus17[31];
assign
s_logisimBus5[49]
=
s_logisimBus17[31];
assign
s_logisimBus5[50]
=
s_logisimBus17[31];
assign
s_logisimBus5[51]
=
s_logisimBus17[31];
assign
s_logisimBus5[52]
=
s_logisimBus17[31];
assign
s_logisimBus5[53]
=
s_logisimBus17[31];
assign
s_logisimBus5[54]
=
s_logisimBus17[31];
assign
s_logisimBus5[55]
=
s_logisimBus17[31];
assign
s_logisimBus5[56]
=
s_logisimBus17[31];
assign
s_logisimBus5[57]
=
s_logisimBus17[31];
assign
s_logisimBus5[58]
=
s_logisimBus17[31];
assign
s_logisimBus5[59]
=
s_logisimBus17[31];
assign
s_logisimBus5[60]
=
s_logisimBus17[31];
assign
s_logisimBus5[61]
=
s_logisimBus17[31];
assign
s_logisimBus5[62]
=
s_logisimBus17[31];
assign
s_logisimBus5[63]
=
s_logisimBus17[31];
assign
s_logisimBus14[5:0]
=
{2'b00,
4'h1};
assign
s_logisimBus22[31:0]
=
32'h00000001;
assign
s_logisimBus25[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus23[31:0]
=
32'h00000000;
assign
s_logisimBus24[31:0]
=
32'hFFFFFFFF;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_1
(.enable(1'b1),
.muxIn_0(s_logisimBus3[63:0]),
.muxIn_1(s_logisimBus18[63:0]),
.muxOut(s_logisimBus12[63:0]),
.sel(s_logisimBus9[0]));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus23[31:0]),
.muxIn_1(s_logisimBus24[31:0]),
.muxOut(s_logisimBus20[63:32]),
.sel(s_logisimBus10[31]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus12[63:0]),
.muxIn_1(s_logisimBus5[63:0]),
.muxOut(s_logisimBus10[63:0]),
.sel(s_logisimNet4));
Shifter_64_bit
#(.shifterMode(2))
ARITH_4
(.dataA(s_logisimBus5[63:0]),
.result(s_logisimBus21[63:0]),
.shiftAmount(s_logisimBus14[5:0]));
Subtractor
#(.extendedBits(33),
.nrOfBits(32))
ARITH_5
(.borrowIn(1'b0),
.borrowOut(),
.dataA(s_logisimBus9[31:0]),
.dataB(s_logisimBus22[31:0]),
.result(s_logisimBus13[31:0]));
Shifter_64_bit
#(.shifterMode(2))
ARITH_6
(.dataA(s_logisimBus5[63:0]),
.result(s_logisimBus18[63:0]),
.shiftAmount(s_logisimBus9[5:0]));
Shifter_64_bit
#(.shifterMode(2))
ARITH_7
(.dataA(s_logisimBus21[63:0]),
.result(s_logisimBus3[63:0]),
.shiftAmount(s_logisimBus13[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_8
(.aEqualsB(s_logisimNet4),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus25[5:0]));
endmodule