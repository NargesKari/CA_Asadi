/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
ROTATE
**
**
**
*****************************************************************************/
module
ROTATE(
a,
b,
ouuut
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[31:0]
b;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[63:0]
ouuut;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[63:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus1;
wire
[31:0]
s_logisimBus2;
wire
[63:0]
s_logisimBus3;
wire
[31:0]
s_logisimBus4;
wire
[31:0]
s_logisimBus5;
wire
[31:0]
s_logisimBus6;
wire
[63:0]
s_logisimBus7;
wire
[63:0]
s_logisimBus8;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
wiring
is
defined
**
*******************************************************************************/
assign
s_logisimBus1[0]
=
s_logisimBus8[0];
assign
s_logisimBus1[10]
=
s_logisimBus8[10];
assign
s_logisimBus1[11]
=
s_logisimBus8[11];
assign
s_logisimBus1[12]
=
s_logisimBus8[12];
assign
s_logisimBus1[13]
=
s_logisimBus8[13];
assign
s_logisimBus1[14]
=
s_logisimBus8[14];
assign
s_logisimBus1[15]
=
s_logisimBus8[15];
assign
s_logisimBus1[16]
=
s_logisimBus8[16];
assign
s_logisimBus1[17]
=
s_logisimBus8[17];
assign
s_logisimBus1[18]
=
s_logisimBus8[18];
assign
s_logisimBus1[19]
=
s_logisimBus8[19];
assign
s_logisimBus1[1]
=
s_logisimBus8[1];
assign
s_logisimBus1[20]
=
s_logisimBus8[20];
assign
s_logisimBus1[21]
=
s_logisimBus8[21];
assign
s_logisimBus1[22]
=
s_logisimBus8[22];
assign
s_logisimBus1[23]
=
s_logisimBus8[23];
assign
s_logisimBus1[24]
=
s_logisimBus8[24];
assign
s_logisimBus1[25]
=
s_logisimBus8[25];
assign
s_logisimBus1[26]
=
s_logisimBus8[26];
assign
s_logisimBus1[27]
=
s_logisimBus8[27];
assign
s_logisimBus1[28]
=
s_logisimBus8[28];
assign
s_logisimBus1[29]
=
s_logisimBus8[29];
assign
s_logisimBus1[2]
=
s_logisimBus8[2];
assign
s_logisimBus1[30]
=
s_logisimBus8[30];
assign
s_logisimBus1[31]
=
s_logisimBus8[31];
assign
s_logisimBus1[3]
=
s_logisimBus8[3];
assign
s_logisimBus1[4]
=
s_logisimBus8[4];
assign
s_logisimBus1[5]
=
s_logisimBus8[5];
assign
s_logisimBus1[6]
=
s_logisimBus8[6];
assign
s_logisimBus1[7]
=
s_logisimBus8[7];
assign
s_logisimBus1[8]
=
s_logisimBus8[8];
assign
s_logisimBus1[9]
=
s_logisimBus8[9];
assign
s_logisimBus3[0]
=
s_logisimBus1[0];
assign
s_logisimBus3[10]
=
s_logisimBus1[10];
assign
s_logisimBus3[11]
=
s_logisimBus1[11];
assign
s_logisimBus3[12]
=
s_logisimBus1[12];
assign
s_logisimBus3[13]
=
s_logisimBus1[13];
assign
s_logisimBus3[14]
=
s_logisimBus1[14];
assign
s_logisimBus3[15]
=
s_logisimBus1[15];
assign
s_logisimBus3[16]
=
s_logisimBus1[16];
assign
s_logisimBus3[17]
=
s_logisimBus1[17];
assign
s_logisimBus3[18]
=
s_logisimBus1[18];
assign
s_logisimBus3[19]
=
s_logisimBus1[19];
assign
s_logisimBus3[1]
=
s_logisimBus1[1];
assign
s_logisimBus3[20]
=
s_logisimBus1[20];
assign
s_logisimBus3[21]
=
s_logisimBus1[21];
assign
s_logisimBus3[22]
=
s_logisimBus1[22];
assign
s_logisimBus3[23]
=
s_logisimBus1[23];
assign
s_logisimBus3[24]
=
s_logisimBus1[24];
assign
s_logisimBus3[25]
=
s_logisimBus1[25];
assign
s_logisimBus3[26]
=
s_logisimBus1[26];
assign
s_logisimBus3[27]
=
s_logisimBus1[27];
assign
s_logisimBus3[28]
=
s_logisimBus1[28];
assign
s_logisimBus3[29]
=
s_logisimBus1[29];
assign
s_logisimBus3[2]
=
s_logisimBus1[2];
assign
s_logisimBus3[30]
=
s_logisimBus1[30];
assign
s_logisimBus3[31]
=
s_logisimBus1[31];
assign
s_logisimBus3[3]
=
s_logisimBus1[3];
assign
s_logisimBus3[4]
=
s_logisimBus1[4];
assign
s_logisimBus3[5]
=
s_logisimBus1[5];
assign
s_logisimBus3[6]
=
s_logisimBus1[6];
assign
s_logisimBus3[7]
=
s_logisimBus1[7];
assign
s_logisimBus3[8]
=
s_logisimBus1[8];
assign
s_logisimBus3[9]
=
s_logisimBus1[9];
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus4[31:0]
=
a;
assign
s_logisimBus5[31:0]
=
b;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
ouuut
=
s_logisimBus3[63:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus6[31:0]
=
32'h00000020;
assign
s_logisimBus3[63:32]
=
32'h00000000;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE_BUS
#(.BubblesMask(2'b00),
.NrOfBits(64))
GATES_1
(.input1(s_logisimBus7[63:0]),
.input2(s_logisimBus0[63:0]),
.result(s_logisimBus8[63:0]));
Subtractor
#(.extendedBits(33),
.nrOfBits(32))
ARITH_2
(.borrowIn(1'b0),
.borrowOut(),
.dataA(s_logisimBus6[31:0]),
.dataB(s_logisimBus5[31:0]),
.result(s_logisimBus2[31:0]));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
SRL2
SRL2_1
(.a(s_logisimBus4[31:0]),
.b(s_logisimBus5[31:0]),
.output1(s_logisimBus7[63:0]));
SLL1
SLL1_1
(.a(s_logisimBus4[31:0]),
.b(s_logisimBus2[31:0]),
.output1(s_logisimBus0[63:0]));
endmodule