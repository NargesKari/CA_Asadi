/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
ALU
**
**
**
*****************************************************************************/
module
ALU(
a,
aluop,
b,
clk,
done,
output_inc,
output_inverted,
res_high,
res_low,
rst
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[3:0]
aluop;
input
[31:0]
b;
input
clk;
input
output_inc;
input
output_inverted;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
done;
output
[31:0]
res_high;
output
[31:0]
res_low;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus1;
wire
[31:0]
s_logisimBus10;
wire
[63:0]
s_logisimBus12;
wire
[63:0]
s_logisimBus14;
wire
[63:0]
s_logisimBus16;
wire
[63:0]
s_logisimBus17;
wire
[63:0]
s_logisimBus18;
wire
[31:0]
s_logisimBus19;
wire
[63:0]
s_logisimBus23;
wire
[63:0]
s_logisimBus24;
wire
[63:0]
s_logisimBus27;
wire
[63:0]
s_logisimBus28;
wire
[3:0]
s_logisimBus30;
wire
[63:0]
s_logisimBus31;
wire
[31:0]
s_logisimBus32;
wire
[63:0]
s_logisimBus33;
wire
[63:0]
s_logisimBus34;
wire
[63:0]
s_logisimBus36;
wire
[63:0]
s_logisimBus37;
wire
[63:0]
s_logisimBus38;
wire
[31:0]
s_logisimBus39;
wire
[31:0]
s_logisimBus40;
wire
[63:0]
s_logisimBus41;
wire
[31:0]
s_logisimBus42;
wire
[63:0]
s_logisimBus44;
wire
[63:0]
s_logisimBus8;
wire
s_logisimNet11;
wire
s_logisimNet21;
wire
s_logisimNet25;
wire
s_logisimNet35;
wire
s_logisimNet43;
wire
s_logisimNet45;
wire
s_logisimNet5;
wire
s_logisimNet6;
wire
s_logisimNet7;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
wiring
is
defined
**
*******************************************************************************/
assign
s_logisimBus14[32]
=
s_logisimBus19[0];
assign
s_logisimBus14[33]
=
s_logisimBus19[1];
assign
s_logisimBus14[34]
=
s_logisimBus19[2];
assign
s_logisimBus14[35]
=
s_logisimBus19[3];
assign
s_logisimBus14[36]
=
s_logisimBus19[4];
assign
s_logisimBus14[37]
=
s_logisimBus19[5];
assign
s_logisimBus14[38]
=
s_logisimBus19[6];
assign
s_logisimBus14[39]
=
s_logisimBus19[7];
assign
s_logisimBus14[40]
=
s_logisimBus19[8];
assign
s_logisimBus14[41]
=
s_logisimBus19[9];
assign
s_logisimBus14[42]
=
s_logisimBus19[10];
assign
s_logisimBus14[43]
=
s_logisimBus19[11];
assign
s_logisimBus14[44]
=
s_logisimBus19[12];
assign
s_logisimBus14[45]
=
s_logisimBus19[13];
assign
s_logisimBus14[46]
=
s_logisimBus19[14];
assign
s_logisimBus14[47]
=
s_logisimBus19[15];
assign
s_logisimBus14[48]
=
s_logisimBus19[16];
assign
s_logisimBus14[49]
=
s_logisimBus19[17];
assign
s_logisimBus14[50]
=
s_logisimBus19[18];
assign
s_logisimBus14[51]
=
s_logisimBus19[19];
assign
s_logisimBus14[52]
=
s_logisimBus19[20];
assign
s_logisimBus14[53]
=
s_logisimBus19[21];
assign
s_logisimBus14[54]
=
s_logisimBus19[22];
assign
s_logisimBus14[55]
=
s_logisimBus19[23];
assign
s_logisimBus14[56]
=
s_logisimBus19[24];
assign
s_logisimBus14[57]
=
s_logisimBus19[25];
assign
s_logisimBus14[58]
=
s_logisimBus19[26];
assign
s_logisimBus14[59]
=
s_logisimBus19[27];
assign
s_logisimBus14[60]
=
s_logisimBus19[28];
assign
s_logisimBus14[61]
=
s_logisimBus19[29];
assign
s_logisimBus14[62]
=
s_logisimBus19[30];
assign
s_logisimBus14[63]
=
s_logisimBus19[31];
assign
s_logisimBus31[32]
=
s_logisimBus19[0];
assign
s_logisimBus31[33]
=
s_logisimBus19[1];
assign
s_logisimBus31[34]
=
s_logisimBus19[2];
assign
s_logisimBus31[35]
=
s_logisimBus19[3];
assign
s_logisimBus31[36]
=
s_logisimBus19[4];
assign
s_logisimBus31[37]
=
s_logisimBus19[5];
assign
s_logisimBus31[38]
=
s_logisimBus19[6];
assign
s_logisimBus31[39]
=
s_logisimBus19[7];
assign
s_logisimBus31[40]
=
s_logisimBus19[8];
assign
s_logisimBus31[41]
=
s_logisimBus19[9];
assign
s_logisimBus31[42]
=
s_logisimBus19[10];
assign
s_logisimBus31[43]
=
s_logisimBus19[11];
assign
s_logisimBus31[44]
=
s_logisimBus19[12];
assign
s_logisimBus31[45]
=
s_logisimBus19[13];
assign
s_logisimBus31[46]
=
s_logisimBus19[14];
assign
s_logisimBus31[47]
=
s_logisimBus19[15];
assign
s_logisimBus31[48]
=
s_logisimBus19[16];
assign
s_logisimBus31[49]
=
s_logisimBus19[17];
assign
s_logisimBus31[50]
=
s_logisimBus19[18];
assign
s_logisimBus31[51]
=
s_logisimBus19[19];
assign
s_logisimBus31[52]
=
s_logisimBus19[20];
assign
s_logisimBus31[53]
=
s_logisimBus19[21];
assign
s_logisimBus31[54]
=
s_logisimBus19[22];
assign
s_logisimBus31[55]
=
s_logisimBus19[23];
assign
s_logisimBus31[56]
=
s_logisimBus19[24];
assign
s_logisimBus31[57]
=
s_logisimBus19[25];
assign
s_logisimBus31[58]
=
s_logisimBus19[26];
assign
s_logisimBus31[59]
=
s_logisimBus19[27];
assign
s_logisimBus31[60]
=
s_logisimBus19[28];
assign
s_logisimBus31[61]
=
s_logisimBus19[29];
assign
s_logisimBus31[62]
=
s_logisimBus19[30];
assign
s_logisimBus31[63]
=
s_logisimBus19[31];
assign
s_logisimBus41[32]
=
s_logisimBus19[0];
assign
s_logisimBus41[33]
=
s_logisimBus19[1];
assign
s_logisimBus41[34]
=
s_logisimBus19[2];
assign
s_logisimBus41[35]
=
s_logisimBus19[3];
assign
s_logisimBus41[36]
=
s_logisimBus19[4];
assign
s_logisimBus41[37]
=
s_logisimBus19[5];
assign
s_logisimBus41[38]
=
s_logisimBus19[6];
assign
s_logisimBus41[39]
=
s_logisimBus19[7];
assign
s_logisimBus41[40]
=
s_logisimBus19[8];
assign
s_logisimBus41[41]
=
s_logisimBus19[9];
assign
s_logisimBus41[42]
=
s_logisimBus19[10];
assign
s_logisimBus41[43]
=
s_logisimBus19[11];
assign
s_logisimBus41[44]
=
s_logisimBus19[12];
assign
s_logisimBus41[45]
=
s_logisimBus19[13];
assign
s_logisimBus41[46]
=
s_logisimBus19[14];
assign
s_logisimBus41[47]
=
s_logisimBus19[15];
assign
s_logisimBus41[48]
=
s_logisimBus19[16];
assign
s_logisimBus41[49]
=
s_logisimBus19[17];
assign
s_logisimBus41[50]
=
s_logisimBus19[18];
assign
s_logisimBus41[51]
=
s_logisimBus19[19];
assign
s_logisimBus41[52]
=
s_logisimBus19[20];
assign
s_logisimBus41[53]
=
s_logisimBus19[21];
assign
s_logisimBus41[54]
=
s_logisimBus19[22];
assign
s_logisimBus41[55]
=
s_logisimBus19[23];
assign
s_logisimBus41[56]
=
s_logisimBus19[24];
assign
s_logisimBus41[57]
=
s_logisimBus19[25];
assign
s_logisimBus41[58]
=
s_logisimBus19[26];
assign
s_logisimBus41[59]
=
s_logisimBus19[27];
assign
s_logisimBus41[60]
=
s_logisimBus19[28];
assign
s_logisimBus41[61]
=
s_logisimBus19[29];
assign
s_logisimBus41[62]
=
s_logisimBus19[30];
assign
s_logisimBus41[63]
=
s_logisimBus19[31];
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus30[3:0]
=
aluop;
assign
s_logisimBus39[31:0]
=
b;
assign
s_logisimBus42[31:0]
=
a;
assign
s_logisimNet25
=
output_inverted;
assign
s_logisimNet35
=
rst;
assign
s_logisimNet43
=
clk;
assign
s_logisimNet45
=
output_inc;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
done
=
s_logisimNet6;
assign
res_high
=
s_logisimBus8[63:32];
assign
res_low
=
s_logisimBus8[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimNet5
=
1'b1;
assign
s_logisimBus19[31:0]
=
32'h00000000;
assign
s_logisimNet11
=
1'b0;
assign
s_logisimBus32[31:0]
=
32'hFFFFFFFF;
assign
s_logisimBus18[63:33]
=
{3'b000,
28'h0000000};
assign
s_logisimBus10[31:0]
=
32'h00000000;
assign
s_logisimBus44[63:0]
=
64'h0000000000000000;
assign
s_logisimBus40
=
~s_logisimBus39;
assign
s_logisimBus34
=
~s_logisimBus23;
assign
s_logisimBus1
=
~s_logisimBus42;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE_BUS
#(.BubblesMask(2'b00),
.NrOfBits(32))
GATES_1
(.input1(s_logisimBus42[31:0]),
.input2(s_logisimBus39[31:0]),
.result(s_logisimBus31[31:0]));
XOR_GATE_BUS_ONEHOT
#(.BubblesMask(2'b00),
.NrOfBits(32))
GATES_2
(.input1(s_logisimBus42[31:0]),
.input2(s_logisimBus39[31:0]),
.result(s_logisimBus14[31:0]));
AND_GATE_BUS
#(.BubblesMask(2'b00),
.NrOfBits(32))
GATES_3
(.input1(s_logisimBus42[31:0]),
.input2(s_logisimBus39[31:0]),
.result(s_logisimBus41[31:0]));
Multiplexer_bus_16
#(.nrOfBits(64))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus18[63:0]),
.muxIn_1(s_logisimBus38[63:0]),
.muxIn_10(s_logisimBus24[63:0]),
.muxIn_11(s_logisimBus16[63:0]),
.muxIn_12(s_logisimBus12[63:0]),
.muxIn_13(64'd0),
.muxIn_14(64'd0),
.muxIn_15(64'd0),
.muxIn_2(s_logisimBus33[63:0]),
.muxIn_3(s_logisimBus36[63:0]),
.muxIn_4(s_logisimBus41[63:0]),
.muxIn_5(s_logisimBus31[63:0]),
.muxIn_6(s_logisimBus14[63:0]),
.muxIn_7(s_logisimBus37[63:0]),
.muxIn_8(s_logisimBus27[63:0]),
.muxIn_9(s_logisimBus28[63:0]),
.muxOut(s_logisimBus23[63:0]),
.sel(s_logisimBus30[3:0]));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus32[31:0]),
.muxIn_1(s_logisimBus10[31:0]),
.muxOut(s_logisimBus38[63:32]),
.sel(s_logisimNet7));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus23[63:0]),
.muxIn_1(s_logisimBus34[63:0]),
.muxOut(s_logisimBus17[63:0]),
.sel(s_logisimNet25));
Adder
#(.extendedBits(65),
.nrOfBits(64))
ARITH_7
(.carryIn(s_logisimNet45),
.carryOut(),
.dataA(s_logisimBus44[63:0]),
.dataB(s_logisimBus17[63:0]),
.result(s_logisimBus8[63:0]));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
mul11
mul11_1
(.a(s_logisimBus42[31:0]),
.b(s_logisimBus39[31:0]),
.mul_out(s_logisimBus33[63:0]));
clooo
clooo_1
(.A(s_logisimBus42[31:0]),
.OUTTTT(s_logisimBus37[63:0]));
clooo
clooo_2
(.A(s_logisimBus1[31:0]),
.OUTTTT(s_logisimBus27[63:0]));
divi
divi_1
(.clk(s_logisimNet43),
.dividend(s_logisimBus42[31:0]),
.divisor(s_logisimBus39[31:0]),
.done(s_logisimNet6),
.quotient(s_logisimBus36[31:0]),
.remainder(s_logisimBus36[63:32]));
ROTATE
ROTATE_1
(.a(s_logisimBus42[31:0]),
.b(s_logisimBus39[31:0]),
.ouuut(s_logisimBus12[63:0]));
CSA
CSA_1
(.A(s_logisimBus42[31:0]),
.B(s_logisimBus39[31:0]),
.SUM(s_logisimBus18[31:0]),
.cin(s_logisimNet11),
.cout(s_logisimBus18[32]));
CSA
CSA_2
(.A(s_logisimBus42[31:0]),
.B(s_logisimBus40[31:0]),
.SUM(s_logisimBus38[31:0]),
.cin(s_logisimNet5),
.cout(s_logisimNet7));
SRA11
SRA11_1
(.a(s_logisimBus42[31:0]),
.b(s_logisimBus39[31:0]),
.output1(s_logisimBus16[63:0]));
SRL2
SRL2_1
(.a(s_logisimBus42[31:0]),
.b(s_logisimBus39[31:0]),
.output1(s_logisimBus24[63:0]));
SLL1
SLL1_1
(.a(s_logisimBus42[31:0]),
.b(s_logisimBus39[31:0]),
.output1(s_logisimBus28[63:0]));
endmodule