/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
PCU
**
**
**
*****************************************************************************/
module
PCU(
ALUOp,
ALUSrc,
Branch,
INS,
Jump,
MemRead,
MemWrite,
MemtoReg,
RegDst,
RegWrite,
clk,
full5,
imm_16,
imm_16_forPC,
isDiv,
isJal,
isMfhi,
isMflo,
isNe,
isRJ,
isSll_shmt,
isSlti,
rd_w,
rs,
rst,
rt,
rt_w,
shamt
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
INS;
input
clk;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[3:0]
ALUOp;
output
ALUSrc;
output
Branch;
output
Jump;
output
MemRead;
output
MemWrite;
output
MemtoReg;
output
RegDst;
output
RegWrite;
output
full5;
output
[15:0]
imm_16;
output
[15:0]
imm_16_forPC;
output
isDiv;
output
isJal;
output
isMfhi;
output
isMflo;
output
isNe;
output
isRJ;
output
isSll_shmt;
output
isSlti;
output
[4:0]
rd_w;
output
[4:0]
rs;
output
[4:0]
rt;
output
[4:0]
rt_w;
output
[4:0]
shamt;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[32:0]
s_logisimBus10;
wire
[32:0]
s_logisimBus11;
wire
[32:0]
s_logisimBus24;
wire
[32:0]
s_logisimBus3;
wire
[32:0]
s_logisimBus4;
wire
[3:0]
s_logisimBus41;
wire
[32:0]
s_logisimBus46;
wire
s_logisimNet0;
wire
s_logisimNet12;
wire
s_logisimNet13;
wire
s_logisimNet16;
wire
s_logisimNet18;
wire
s_logisimNet25;
wire
s_logisimNet27;
wire
s_logisimNet28;
wire
s_logisimNet29;
wire
s_logisimNet37;
wire
s_logisimNet39;
wire
s_logisimNet40;
wire
s_logisimNet45;
wire
s_logisimNet47;
wire
s_logisimNet48;
wire
s_logisimNet49;
wire
s_logisimNet50;
wire
s_logisimNet51;
wire
s_logisimNet52;
wire
s_logisimNet54;
wire
s_logisimNet55;
wire
s_logisimNet56;
wire
s_logisimNet57;
wire
s_logisimNet58;
wire
s_logisimNet6;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus24[31:0]
=
INS;
assign
s_logisimNet0
=
clk;
assign
s_logisimNet6
=
rst;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
ALUOp
=
s_logisimBus41[3:0];
assign
ALUSrc
=
s_logisimNet12;
assign
Branch
=
s_logisimNet47;
assign
Jump
=
s_logisimNet28;
assign
MemRead
=
s_logisimNet51;
assign
MemWrite
=
s_logisimNet27;
assign
MemtoReg
=
s_logisimNet39;
assign
RegDst
=
s_logisimNet45;
assign
RegWrite
=
s_logisimNet54;
assign
full5
=
s_logisimBus46[32];
assign
imm_16
=
s_logisimBus3[15:0];
assign
imm_16_forPC
=
s_logisimBus11[15:0];
assign
isDiv
=
s_logisimNet13;
assign
isJal
=
s_logisimNet40;
assign
isMfhi
=
s_logisimNet55;
assign
isMflo
=
s_logisimNet56;
assign
isNe
=
s_logisimNet48;
assign
isRJ
=
s_logisimNet52;
assign
isSll_shmt
=
s_logisimNet37;
assign
isSlti
=
s_logisimNet29;
assign
rd_w
=
s_logisimBus10[15:11];
assign
rs
=
s_logisimBus4[25:21];
assign
rt
=
s_logisimBus4[20:16];
assign
rt_w
=
s_logisimBus10[20:16];
assign
shamt
=
s_logisimBus3[10:6];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimNet49
=
1'b1;
assign
s_logisimNet58
=
1'b1;
assign
s_logisimNet25
=
1'b1;
assign
s_logisimBus24[32]
=
1'b1;
assign
s_logisimNet18
=
1'b1;
assign
s_logisimNet16
=
1'b1;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(33))
ALU
(.clock(s_logisimNet0),
.clockEnable(s_logisimNet49),
.d(s_logisimBus3[32:0]),
.q(s_logisimBus11[32:0]),
.reset(s_logisimNet6),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(33))
D_MEM
(.clock(s_logisimNet0),
.clockEnable(s_logisimNet58),
.d(s_logisimBus11[32:0]),
.q(s_logisimBus10[32:0]),
.reset(s_logisimNet6),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(33))
RW
(.clock(s_logisimNet0),
.clockEnable(s_logisimNet25),
.d(s_logisimBus10[32:0]),
.q(s_logisimBus46[32:0]),
.reset(s_logisimNet6),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(33))
I_MEM
(.clock(s_logisimNet0),
.clockEnable(s_logisimNet18),
.d(s_logisimBus24[32:0]),
.q(s_logisimBus4[32:0]),
.reset(s_logisimNet6),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(33))
REGS
(.clock(s_logisimNet0),
.clockEnable(s_logisimNet16),
.d(s_logisimBus4[32:0]),
.q(s_logisimBus3[32:0]),
.reset(s_logisimNet6),
.tick(1'b1));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
CU
CU_2
(.ALUSrc(s_logisimNet12),
.AlUOp(s_logisimBus41[3:0]),
.Branch(),
.IsNe(),
.Jump(),
.MemRead(),
.MemWrite(),
.MemtoReg(),
.RegDst(),
.RegWrite(),
.func(s_logisimBus3[5:0]),
.isDiv(s_logisimNet13),
.isJal(),
.isMfhi(),
.isMflo(),
.isRJ(),
.isSll_shmt(s_logisimNet37),
.isSlti(),
.op_code(s_logisimBus3[31:26]));
CU
CU_3
(.ALUSrc(),
.AlUOp(),
.Branch(s_logisimNet47),
.IsNe(s_logisimNet48),
.Jump(s_logisimNet28),
.MemRead(s_logisimNet51),
.MemWrite(s_logisimNet27),
.MemtoReg(),
.RegDst(),
.RegWrite(),
.func(s_logisimBus11[5:0]),
.isDiv(),
.isJal(),
.isMfhi(),
.isMflo(),
.isRJ(s_logisimNet52),
.isSll_shmt(),
.isSlti(),
.op_code(s_logisimBus11[31:26]));
CU
CU_4
(.ALUSrc(),
.AlUOp(),
.Branch(),
.IsNe(),
.Jump(),
.MemRead(),
.MemWrite(),
.MemtoReg(s_logisimNet39),
.RegDst(s_logisimNet45),
.RegWrite(s_logisimNet54),
.func(s_logisimBus10[5:0]),
.isDiv(),
.isJal(s_logisimNet40),
.isMfhi(s_logisimNet55),
.isMflo(s_logisimNet56),
.isRJ(),
.isSll_shmt(),
.isSlti(s_logisimNet29),
.op_code(s_logisimBus10[31:26]));
CU
CU_5
(.ALUSrc(),
.AlUOp(),
.Branch(),
.IsNe(),
.Jump(),
.MemRead(),
.MemWrite(),
.MemtoReg(),
.RegDst(),
.RegWrite(),
.func(s_logisimBus46[5:0]),
.isDiv(),
.isJal(),
.isMfhi(),
.isMflo(),
.isRJ(),
.isSll_shmt(),
.isSlti(),
.op_code(s_logisimBus46[31:26]));
CU
CU_1
(.ALUSrc(),
.AlUOp(),
.Branch(),
.IsNe(),
.Jump(),
.MemRead(),
.MemWrite(),
.MemtoReg(),
.RegDst(),
.RegWrite(),
.func(s_logisimBus4[5:0]),
.isDiv(),
.isJal(),
.isMfhi(),
.isMflo(),
.isRJ(),
.isSll_shmt(),
.isSlti(),
.op_code(s_logisimBus4[31:26]));
endmodule