/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
PC_Update
**
**
**
*****************************************************************************/
module
PC_Update(
Branch,
Eq,
Imm,
Jump,
PC,
PC_out,
clk,
divIsActive,
isNe
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
Branch;
input
[31:0]
Eq;
input
[15:0]
Imm;
input
Jump;
input
[8:0]
PC;
input
clk;
input
divIsActive;
input
isNe;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[8:0]
PC_out;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[15:0]
s_logisimBus0;
wire
[8:0]
s_logisimBus1;
wire
[8:0]
s_logisimBus12;
wire
[8:0]
s_logisimBus15;
wire
[31:0]
s_logisimBus16;
wire
[8:0]
s_logisimBus17;
wire
[8:0]
s_logisimBus19;
wire
[8:0]
s_logisimBus2;
wire
[8:0]
s_logisimBus20;
wire
[31:0]
s_logisimBus24;
wire
[8:0]
s_logisimBus4;
wire
[8:0]
s_logisimBus6;
wire
[8:0]
s_logisimBus7;
wire
[8:0]
s_logisimBus8;
wire
[8:0]
s_logisimBus9;
wire
s_logisimNet10;
wire
s_logisimNet11;
wire
s_logisimNet13;
wire
s_logisimNet14;
wire
s_logisimNet18;
wire
s_logisimNet21;
wire
s_logisimNet22;
wire
s_logisimNet23;
wire
s_logisimNet25;
wire
s_logisimNet3;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus0[15:0]
=
Imm;
assign
s_logisimBus16[31:0]
=
Eq;
assign
s_logisimBus2[8:0]
=
PC;
assign
s_logisimNet10
=
Branch;
assign
s_logisimNet11
=
Jump;
assign
s_logisimNet14
=
isNe;
assign
s_logisimNet25
=
clk;
assign
s_logisimNet3
=
divIsActive;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
PC_out
=
s_logisimBus17[8:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus20[8:0]
=
{1'b0,
8'h01};
assign
s_logisimNet22
=
1'b0;
assign
s_logisimBus24[31:0]
=
32'h00000000;
assign
s_logisimNet23
=
1'b0;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
XOR_GATE_ONEHOT
#(.BubblesMask(2'b00))
GATES_1
(.input1(s_logisimNet14),
.input2(s_logisimNet13),
.result(s_logisimNet21));
AND_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet10),
.input2(s_logisimNet21),
.result(s_logisimNet18));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus1[8:0]),
.muxIn_1(s_logisimBus12[8:0]),
.muxOut(s_logisimBus7[8:0]),
.sel(s_logisimNet18));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus7[8:0]),
.muxIn_1(s_logisimBus0[8:0]),
.muxOut(s_logisimBus19[8:0]),
.sel(s_logisimNet11));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus19[8:0]),
.muxIn_1(s_logisimBus2[8:0]),
.muxOut(s_logisimBus17[8:0]),
.sel(s_logisimNet3));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_6
(.carryIn(s_logisimNet22),
.carryOut(),
.dataA(s_logisimBus20[8:0]),
.dataB(s_logisimBus2[8:0]),
.result(s_logisimBus1[8:0]));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_7
(.carryIn(s_logisimNet23),
.carryOut(),
.dataA(s_logisimBus15[8:0]),
.dataB(s_logisimBus0[8:0]),
.result(s_logisimBus12[8:0]));
Comparator
#(.nrOfBits(32),
.twosComplement(1))
ARITH_8
(.aEqualsB(s_logisimNet13),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus16[31:0]),
.dataB(s_logisimBus24[31:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
MEMORY_9
(.clock(s_logisimNet25),
.clockEnable(1'b1),
.d(s_logisimBus1[8:0]),
.q(s_logisimBus6[8:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
MEMORY_10
(.clock(s_logisimNet25),
.clockEnable(1'b1),
.d(s_logisimBus6[8:0]),
.q(s_logisimBus8[8:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
MEMORY_11
(.clock(s_logisimNet25),
.clockEnable(1'b1),
.d(s_logisimBus8[8:0]),
.q(s_logisimBus9[8:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
MEMORY_12
(.clock(s_logisimNet25),
.clockEnable(1'b1),
.d(s_logisimBus9[8:0]),
.q(s_logisimBus4[8:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
MEMORY_13
(.clock(s_logisimNet25),
.clockEnable(1'b1),
.d(s_logisimBus4[8:0]),
.q(s_logisimBus15[8:0]),
.reset(1'b0),
.tick(1'b1));
endmodule