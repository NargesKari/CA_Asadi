/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
main
**
**
**
*****************************************************************************/
module
main(
InstDone,
Jen,
Jin,
Jout,
R1,
R10,
R11,
R12,
R13,
R14,
R15,
R16,
R17,
R18,
R19,
R2,
R20,
R21,
R22,
R23,
R24,
R25,
R26,
R27,
R28,
R29,
R3,
R30,
R31,
R4,
R5,
R6,
R7,
R8,
R9,
clk,
rst
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
Jen;
input
[31:0]
Jin;
input
clk;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
InstDone;
output
[31:0]
Jout;
output
[31:0]
R1;
output
[31:0]
R10;
output
[31:0]
R11;
output
[31:0]
R12;
output
[31:0]
R13;
output
[31:0]
R14;
output
[31:0]
R15;
output
[31:0]
R16;
output
[31:0]
R17;
output
[31:0]
R18;
output
[31:0]
R19;
output
[31:0]
R2;
output
[31:0]
R20;
output
[31:0]
R21;
output
[31:0]
R22;
output
[31:0]
R23;
output
[31:0]
R24;
output
[31:0]
R25;
output
[31:0]
R26;
output
[31:0]
R27;
output
[31:0]
R28;
output
[31:0]
R29;
output
[31:0]
R3;
output
[31:0]
R30;
output
[31:0]
R31;
output
[31:0]
R4;
output
[31:0]
R5;
output
[31:0]
R6;
output
[31:0]
R7;
output
[31:0]
R8;
output
[31:0]
R9;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus1;
wire
[31:0]
s_logisimBus10;
wire
[31:0]
s_logisimBus100;
wire
[3:0]
s_logisimBus101;
wire
[5:0]
s_logisimBus102;
wire
[4:0]
s_logisimBus103;
wire
[31:0]
s_logisimBus11;
wire
[31:0]
s_logisimBus12;
wire
[31:0]
s_logisimBus13;
wire
[31:0]
s_logisimBus14;
wire
[31:0]
s_logisimBus15;
wire
[31:0]
s_logisimBus16;
wire
[31:0]
s_logisimBus17;
wire
[31:0]
s_logisimBus18;
wire
[31:0]
s_logisimBus19;
wire
[31:0]
s_logisimBus20;
wire
[31:0]
s_logisimBus21;
wire
[31:0]
s_logisimBus22;
wire
[15:0]
s_logisimBus23;
wire
[4:0]
s_logisimBus24;
wire
[4:0]
s_logisimBus25;
wire
[8:0]
s_logisimBus26;
wire
[15:0]
s_logisimBus28;
wire
[31:0]
s_logisimBus3;
wire
[31:0]
s_logisimBus31;
wire
[31:0]
s_logisimBus32;
wire
[4:0]
s_logisimBus33;
wire
[31:0]
s_logisimBus34;
wire
[5:0]
s_logisimBus38;
wire
[31:0]
s_logisimBus4;
wire
[31:0]
s_logisimBus41;
wire
[31:0]
s_logisimBus42;
wire
[31:0]
s_logisimBus44;
wire
[31:0]
s_logisimBus46;
wire
[31:0]
s_logisimBus49;
wire
[31:0]
s_logisimBus5;
wire
[31:0]
s_logisimBus51;
wire
[31:0]
s_logisimBus52;
wire
[31:0]
s_logisimBus53;
wire
[31:0]
s_logisimBus54;
wire
[31:0]
s_logisimBus55;
wire
[31:0]
s_logisimBus56;
wire
[31:0]
s_logisimBus57;
wire
[31:0]
s_logisimBus58;
wire
[31:0]
s_logisimBus59;
wire
[31:0]
s_logisimBus6;
wire
[31:0]
s_logisimBus60;
wire
[31:0]
s_logisimBus61;
wire
[31:0]
s_logisimBus62;
wire
[31:0]
s_logisimBus63;
wire
[31:0]
s_logisimBus64;
wire
[31:0]
s_logisimBus65;
wire
[31:0]
s_logisimBus66;
wire
[31:0]
s_logisimBus67;
wire
[4:0]
s_logisimBus68;
wire
[4:0]
s_logisimBus69;
wire
[31:0]
s_logisimBus7;
wire
[31:0]
s_logisimBus72;
wire
[4:0]
s_logisimBus76;
wire
[31:0]
s_logisimBus8;
wire
[31:0]
s_logisimBus80;
wire
[31:0]
s_logisimBus82;
wire
[31:0]
s_logisimBus85;
wire
[31:0]
s_logisimBus86;
wire
[31:0]
s_logisimBus88;
wire
[31:0]
s_logisimBus9;
wire
[31:0]
s_logisimBus90;
wire
[31:0]
s_logisimBus91;
wire
[4:0]
s_logisimBus97;
wire
[4:0]
s_logisimBus98;
wire
[31:0]
s_logisimBus99;
wire
s_logisimNet104;
wire
s_logisimNet2;
wire
s_logisimNet27;
wire
s_logisimNet29;
wire
s_logisimNet30;
wire
s_logisimNet35;
wire
s_logisimNet36;
wire
s_logisimNet37;
wire
s_logisimNet39;
wire
s_logisimNet43;
wire
s_logisimNet45;
wire
s_logisimNet48;
wire
s_logisimNet50;
wire
s_logisimNet71;
wire
s_logisimNet73;
wire
s_logisimNet74;
wire
s_logisimNet75;
wire
s_logisimNet77;
wire
s_logisimNet78;
wire
s_logisimNet79;
wire
s_logisimNet81;
wire
s_logisimNet83;
wire
s_logisimNet87;
wire
s_logisimNet89;
wire
s_logisimNet92;
wire
s_logisimNet93;
wire
s_logisimNet94;
wire
s_logisimNet95;
wire
s_logisimNet96;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus1[31:0]
=
Jin;
assign
s_logisimNet104
=
clk;
assign
s_logisimNet37
=
Jen;
assign
s_logisimNet96
=
rst;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
InstDone
=
s_logisimNet78;
assign
Jout
=
s_logisimBus5[31:0];
assign
R1
=
s_logisimBus53[31:0];
assign
R10
=
s_logisimBus10[31:0];
assign
R11
=
s_logisimBus57[31:0];
assign
R12
=
s_logisimBus11[31:0];
assign
R13
=
s_logisimBus58[31:0];
assign
R14
=
s_logisimBus12[31:0];
assign
R15
=
s_logisimBus59[31:0];
assign
R16
=
s_logisimBus13[31:0];
assign
R17
=
s_logisimBus60[31:0];
assign
R18
=
s_logisimBus14[31:0];
assign
R19
=
s_logisimBus61[31:0];
assign
R2
=
s_logisimBus8[31:0];
assign
R20
=
s_logisimBus15[31:0];
assign
R21
=
s_logisimBus62[31:0];
assign
R22
=
s_logisimBus16[31:0];
assign
R23
=
s_logisimBus63[31:0];
assign
R24
=
s_logisimBus17[31:0];
assign
R25
=
s_logisimBus64[31:0];
assign
R26
=
s_logisimBus18[31:0];
assign
R27
=
s_logisimBus65[31:0];
assign
R28
=
s_logisimBus19[31:0];
assign
R29
=
s_logisimBus66[31:0];
assign
R3
=
s_logisimBus54[31:0];
assign
R30
=
s_logisimBus20[31:0];
assign
R31
=
s_logisimBus67[31:0];
assign
R4
=
s_logisimBus7[31:0];
assign
R5
=
s_logisimBus55[31:0];
assign
R6
=
s_logisimBus9[31:0];
assign
R7
=
s_logisimBus52[31:0];
assign
R8
=
s_logisimBus6[31:0];
assign
R9
=
s_logisimBus56[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus76[4:0]
=
{1'b1,
4'hF};
assign
s_logisimBus91[31:0]
=
32'h00000000;
assign
s_logisimBus68[4:0]
=
{1'b0,
4'h0};
assign
s_logisimBus42[0]
=
s_logisimNet35;
assign
s_logisimBus42[1]
=
1'b0;
assign
s_logisimBus42[2]
=
1'b0;
assign
s_logisimBus42[3]
=
1'b0;
assign
s_logisimBus42[4]
=
1'b0;
assign
s_logisimBus42[5]
=
1'b0;
assign
s_logisimBus42[6]
=
1'b0;
assign
s_logisimBus42[7]
=
1'b0;
assign
s_logisimBus42[8]
=
1'b0;
assign
s_logisimBus42[9]
=
1'b0;
assign
s_logisimBus42[10]
=
1'b0;
assign
s_logisimBus42[11]
=
1'b0;
assign
s_logisimBus42[12]
=
1'b0;
assign
s_logisimBus42[13]
=
1'b0;
assign
s_logisimBus42[14]
=
1'b0;
assign
s_logisimBus42[15]
=
1'b0;
assign
s_logisimBus42[16]
=
1'b0;
assign
s_logisimBus42[17]
=
1'b0;
assign
s_logisimBus42[18]
=
1'b0;
assign
s_logisimBus42[19]
=
1'b0;
assign
s_logisimBus42[20]
=
1'b0;
assign
s_logisimBus42[21]
=
1'b0;
assign
s_logisimBus42[22]
=
1'b0;
assign
s_logisimBus42[23]
=
1'b0;
assign
s_logisimBus42[24]
=
1'b0;
assign
s_logisimBus42[25]
=
1'b0;
assign
s_logisimBus42[26]
=
1'b0;
assign
s_logisimBus42[27]
=
1'b0;
assign
s_logisimBus42[28]
=
1'b0;
assign
s_logisimBus42[29]
=
1'b0;
assign
s_logisimBus42[30]
=
1'b0;
assign
s_logisimBus42[31]
=
1'b0;
assign
s_logisimBus90[31:9]
=
{3'b000,
20'h00000};
assign
s_logisimNet92
=
1'b1;
assign
s_logisimBus82[31:0]
=
32'h00000000;
assign
s_logisimNet2
=
1'b1;
assign
s_logisimBus85[0]
=
s_logisimBus23[0];
assign
s_logisimBus85[1]
=
s_logisimBus23[1];
assign
s_logisimBus85[2]
=
s_logisimBus23[2];
assign
s_logisimBus85[3]
=
s_logisimBus23[3];
assign
s_logisimBus85[4]
=
s_logisimBus23[4];
assign
s_logisimBus85[5]
=
s_logisimBus23[5];
assign
s_logisimBus85[6]
=
s_logisimBus23[6];
assign
s_logisimBus85[7]
=
s_logisimBus23[7];
assign
s_logisimBus85[8]
=
s_logisimBus23[8];
assign
s_logisimBus85[9]
=
s_logisimBus23[9];
assign
s_logisimBus85[10]
=
s_logisimBus23[10];
assign
s_logisimBus85[11]
=
s_logisimBus23[11];
assign
s_logisimBus85[12]
=
s_logisimBus23[12];
assign
s_logisimBus85[13]
=
s_logisimBus23[13];
assign
s_logisimBus85[14]
=
s_logisimBus23[14];
assign
s_logisimBus85[15]
=
s_logisimBus23[15];
assign
s_logisimBus85[16]
=
s_logisimBus23[15];
assign
s_logisimBus85[17]
=
s_logisimBus23[15];
assign
s_logisimBus85[18]
=
s_logisimBus23[15];
assign
s_logisimBus85[19]
=
s_logisimBus23[15];
assign
s_logisimBus85[20]
=
s_logisimBus23[15];
assign
s_logisimBus85[21]
=
s_logisimBus23[15];
assign
s_logisimBus85[22]
=
s_logisimBus23[15];
assign
s_logisimBus85[23]
=
s_logisimBus23[15];
assign
s_logisimBus85[24]
=
s_logisimBus23[15];
assign
s_logisimBus85[25]
=
s_logisimBus23[15];
assign
s_logisimBus85[26]
=
s_logisimBus23[15];
assign
s_logisimBus85[27]
=
s_logisimBus23[15];
assign
s_logisimBus85[28]
=
s_logisimBus23[15];
assign
s_logisimBus85[29]
=
s_logisimBus23[15];
assign
s_logisimBus85[30]
=
s_logisimBus23[15];
assign
s_logisimBus85[31]
=
s_logisimBus23[15];
assign
s_logisimBus72[0]
=
s_logisimBus25[0];
assign
s_logisimBus72[1]
=
s_logisimBus25[1];
assign
s_logisimBus72[2]
=
s_logisimBus25[2];
assign
s_logisimBus72[3]
=
s_logisimBus25[3];
assign
s_logisimBus72[4]
=
s_logisimBus25[4];
assign
s_logisimBus72[5]
=
s_logisimBus25[4];
assign
s_logisimBus72[6]
=
s_logisimBus25[4];
assign
s_logisimBus72[7]
=
s_logisimBus25[4];
assign
s_logisimBus72[8]
=
s_logisimBus25[4];
assign
s_logisimBus72[9]
=
s_logisimBus25[4];
assign
s_logisimBus72[10]
=
s_logisimBus25[4];
assign
s_logisimBus72[11]
=
s_logisimBus25[4];
assign
s_logisimBus72[12]
=
s_logisimBus25[4];
assign
s_logisimBus72[13]
=
s_logisimBus25[4];
assign
s_logisimBus72[14]
=
s_logisimBus25[4];
assign
s_logisimBus72[15]
=
s_logisimBus25[4];
assign
s_logisimBus72[16]
=
s_logisimBus25[4];
assign
s_logisimBus72[17]
=
s_logisimBus25[4];
assign
s_logisimBus72[18]
=
s_logisimBus25[4];
assign
s_logisimBus72[19]
=
s_logisimBus25[4];
assign
s_logisimBus72[20]
=
s_logisimBus25[4];
assign
s_logisimBus72[21]
=
s_logisimBus25[4];
assign
s_logisimBus72[22]
=
s_logisimBus25[4];
assign
s_logisimBus72[23]
=
s_logisimBus25[4];
assign
s_logisimBus72[24]
=
s_logisimBus25[4];
assign
s_logisimBus72[25]
=
s_logisimBus25[4];
assign
s_logisimBus72[26]
=
s_logisimBus25[4];
assign
s_logisimBus72[27]
=
s_logisimBus25[4];
assign
s_logisimBus72[28]
=
s_logisimBus25[4];
assign
s_logisimBus72[29]
=
s_logisimBus25[4];
assign
s_logisimBus72[30]
=
s_logisimBus25[4];
assign
s_logisimBus72[31]
=
s_logisimBus25[4];
assign
s_logisimNet94
=
1'b0;
assign
s_logisimNet95
=
1'b0;
assign
s_logisimNet78
=
~s_logisimNet79;
assign
s_logisimNet87
=
~s_logisimNet74;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE
#(.BubblesMask(2'b00))
GATES_1
(.input1(s_logisimNet87),
.input2(s_logisimNet73),
.result(s_logisimNet79));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus98[4:0]),
.muxIn_1(s_logisimBus103[4:0]),
.muxOut(s_logisimBus33[4:0]),
.sel(s_logisimNet36));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus33[4:0]),
.muxIn_1(s_logisimBus76[4:0]),
.muxOut(s_logisimBus24[4:0]),
.sel(s_logisimNet30));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus68[4:0]),
.muxIn_1(s_logisimBus24[4:0]),
.muxOut(s_logisimBus69[4:0]),
.sel(s_logisimNet89));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus86[31:0]),
.muxIn_1(s_logisimBus32[31:0]),
.muxOut(s_logisimBus0[31:0]),
.sel(s_logisimNet83));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus0[31:0]),
.muxIn_1(s_logisimBus42[31:0]),
.muxOut(s_logisimBus80[31:0]),
.sel(s_logisimNet50));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_7
(.enable(1'b1),
.muxIn_0(s_logisimBus80[31:0]),
.muxIn_1(s_logisimBus88[31:0]),
.muxOut(s_logisimBus3[31:0]),
.sel(s_logisimNet81));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus3[31:0]),
.muxIn_1(s_logisimBus51[31:0]),
.muxOut(s_logisimBus46[31:0]),
.sel(s_logisimNet39));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_9
(.enable(1'b1),
.muxIn_0(s_logisimBus46[31:0]),
.muxIn_1(s_logisimBus21[31:0]),
.muxOut(s_logisimBus4[31:0]),
.sel(s_logisimNet30));
Multiplexer_bus_2
#(.nrOfBits(16))
PLEXERS_10
(.enable(1'b1),
.muxIn_0(s_logisimBus23[15:0]),
.muxIn_1(s_logisimBus99[15:0]),
.muxOut(s_logisimBus28[15:0]),
.sel(s_logisimNet77));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_11
(.enable(1'b1),
.muxIn_0(s_logisimBus100[31:0]),
.muxIn_1(s_logisimBus85[31:0]),
.muxOut(s_logisimBus44[31:0]),
.sel(s_logisimNet27));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_12
(.enable(1'b1),
.muxIn_0(s_logisimBus44[31:0]),
.muxIn_1(s_logisimBus72[31:0]),
.muxOut(s_logisimBus49[31:0]),
.sel(s_logisimNet45));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_13
(.enable(1'b1),
.muxIn_0(s_logisimBus99[31:0]),
.muxIn_1(s_logisimBus100[31:0]),
.muxOut(s_logisimBus22[31:0]),
.sel(s_logisimNet45));
Comparator
#(.nrOfBits(32),
.twosComplement(1))
ARITH_14
(.aEqualsB(),
.aGreaterThanB(s_logisimNet35),
.aLessThanB(),
.dataA(s_logisimBus91[31:0]),
.dataB(s_logisimBus86[31:0]));
Adder
#(.extendedBits(33),
.nrOfBits(32))
ARITH_15
(.carryIn(s_logisimNet2),
.carryOut(),
.dataA(s_logisimBus90[31:0]),
.dataB(s_logisimBus82[31:0]),
.result(s_logisimBus21[31:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
programCounter
(.clock(s_logisimNet104),
.clockEnable(s_logisimNet92),
.d(s_logisimBus26[8:0]),
.q(s_logisimBus90[8:0]),
.reset(s_logisimNet96),
.tick(1'b1));
D_FLIPFLOP
#(.invertClockEnable(0))
MEMORY_17
(.clock(s_logisimNet104),
.d(s_logisimNet93),
.preset(1'b0),
.q(s_logisimNet74),
.qBar(),
.reset(s_logisimNet96),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_18
(.clock(s_logisimNet104),
.clockEnable(s_logisimNet73),
.d(s_logisimBus86[31:0]),
.q(s_logisimBus88[31:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_19
(.clock(s_logisimNet104),
.clockEnable(s_logisimNet73),
.d(s_logisimBus41[31:0]),
.q(s_logisimBus51[31:0]),
.reset(1'b0),
.tick(1'b1));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
ALU
ALU_1
(.a(s_logisimBus22[31:0]),
.aluop(s_logisimBus101[3:0]),
.b(s_logisimBus49[31:0]),
.clk(s_logisimNet104),
.done(s_logisimNet93),
.output_inc(s_logisimNet94),
.output_inverted(s_logisimNet95),
.res_high(s_logisimBus41[31:0]),
.res_low(s_logisimBus86[31:0]),
.rst(s_logisimNet96));
regfile
RF
(.Aread0(s_logisimBus97[4:0]),
.Aread1(s_logisimBus98[4:0]),
.Awrite(s_logisimBus69[4:0]),
.Dread0(s_logisimBus99[31:0]),
.Dread1(s_logisimBus100[31:0]),
.Dwrite(s_logisimBus4[31:0]),
.R1(s_logisimBus53[31:0]),
.R10(s_logisimBus10[31:0]),
.R11(s_logisimBus57[31:0]),
.R12(s_logisimBus11[31:0]),
.R13(s_logisimBus58[31:0]),
.R14(s_logisimBus12[31:0]),
.R15(s_logisimBus59[31:0]),
.R16(s_logisimBus13[31:0]),
.R17(s_logisimBus60[31:0]),
.R18(s_logisimBus14[31:0]),
.R19(s_logisimBus61[31:0]),
.R2(s_logisimBus8[31:0]),
.R20(s_logisimBus15[31:0]),
.R21(s_logisimBus62[31:0]),
.R22(s_logisimBus16[31:0]),
.R23(s_logisimBus63[31:0]),
.R24(s_logisimBus17[31:0]),
.R25(s_logisimBus64[31:0]),
.R26(s_logisimBus18[31:0]),
.R27(s_logisimBus65[31:0]),
.R28(s_logisimBus19[31:0]),
.R29(s_logisimBus66[31:0]),
.R3(s_logisimBus54[31:0]),
.R30(s_logisimBus20[31:0]),
.R31(s_logisimBus67[31:0]),
.R4(s_logisimBus7[31:0]),
.R5(s_logisimBus55[31:0]),
.R6(s_logisimBus9[31:0]),
.R7(s_logisimBus52[31:0]),
.R8(s_logisimBus6[31:0]),
.R9(s_logisimBus56[31:0]),
.clk(s_logisimNet104),
.rst(s_logisimNet96));
CU
Control_Unit
(.ALUSrc(s_logisimNet27),
.AlUOp(s_logisimBus101[3:0]),
.Branch(s_logisimNet48),
.IsNe(s_logisimNet75),
.Jump(s_logisimNet71),
.MemRead(s_logisimNet29),
.MemWrite(s_logisimNet43),
.MemtoReg(s_logisimNet83),
.RegDst(s_logisimNet36),
.RegWrite(s_logisimNet89),
.func(s_logisimBus102[5:0]),
.isDiv(s_logisimNet73),
.isJal(s_logisimNet30),
.isMfhi(s_logisimNet39),
.isMflo(s_logisimNet81),
.isRJ(s_logisimNet77),
.isSll_shmt(s_logisimNet45),
.isSlti(s_logisimNet50),
.op_code(s_logisimBus38[5:0]));
INC_decoder
INC
(.fuunc(s_logisimBus102[5:0]),
.imm(s_logisimBus23[15:0]),
.inc(s_logisimBus34[31:0]),
.op(s_logisimBus38[5:0]),
.rd(s_logisimBus103[4:0]),
.rs(s_logisimBus97[4:0]),
.rt(s_logisimBus98[4:0]),
.shamt(s_logisimBus25[4:0]));
jtag_ram512
I_mem
(.Addr(s_logisimBus90[8:0]),
.Din(32'd0),
.Dout(s_logisimBus34[31:0]),
.Jen(s_logisimNet37),
.Jin(s_logisimBus1[31:0]),
.Jout(s_logisimBus31[31:0]),
.Wen(1'b0),
.clk(s_logisimNet104));
jtag_ram512
D_mem
(.Addr(s_logisimBus86[8:0]),
.Din(s_logisimBus100[31:0]),
.Dout(s_logisimBus32[31:0]),
.Jen(s_logisimNet37),
.Jin(s_logisimBus31[31:0]),
.Jout(s_logisimBus5[31:0]),
.Wen(s_logisimNet43),
.clk(s_logisimNet104));
PC_Update
PC_Update_1
(.Branch(s_logisimNet48),
.Eq(s_logisimBus86[31:0]),
.Imm(s_logisimBus28[15:0]),
.Jump(s_logisimNet71),
.PC(s_logisimBus90[8:0]),
.PC_out(s_logisimBus26[8:0]),
.divIsActive(s_logisimNet79),
.isNe(s_logisimNet75));
endmodule