/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
PC_Update
**
**
**
*****************************************************************************/
module
PC_Update(
Branch,
Eq,
Imm,
Jump,
PC,
PC_out,
divIsActive
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
Branch;
input
[31:0]
Eq;
input
[15:0]
Imm;
input
Jump;
input
[8:0]
PC;
input
divIsActive;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[8:0]
PC_out;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[15:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus11;
wire
[8:0]
s_logisimBus12;
wire
[8:0]
s_logisimBus14;
wire
[8:0]
s_logisimBus15;
wire
[8:0]
s_logisimBus2;
wire
[8:0]
s_logisimBus4;
wire
[8:0]
s_logisimBus5;
wire
[8:0]
s_logisimBus8;
wire
[31:0]
s_logisimBus9;
wire
s_logisimNet10;
wire
s_logisimNet13;
wire
s_logisimNet16;
wire
s_logisimNet17;
wire
s_logisimNet3;
wire
s_logisimNet6;
wire
s_logisimNet7;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus0[15:0]
=
Imm;
assign
s_logisimBus11[31:0]
=
Eq;
assign
s_logisimBus2[8:0]
=
PC;
assign
s_logisimNet3
=
divIsActive;
assign
s_logisimNet6
=
Jump;
assign
s_logisimNet7
=
Branch;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
PC_out
=
s_logisimBus15[8:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus14[8:0]
=
{1'b0,
8'h01};
assign
s_logisimNet16
=
1'b0;
assign
s_logisimNet17
=
1'b0;
assign
s_logisimBus9[31:0]
=
32'h00000000;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE
#(.BubblesMask(2'b10))
GATES_1
(.input1(s_logisimNet7),
.input2(s_logisimNet13),
.result(s_logisimNet10));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus5[8:0]),
.muxIn_1(s_logisimBus8[8:0]),
.muxOut(s_logisimBus4[8:0]),
.sel(s_logisimNet10));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus4[8:0]),
.muxIn_1(s_logisimBus0[8:0]),
.muxOut(s_logisimBus12[8:0]),
.sel(s_logisimNet6));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus12[8:0]),
.muxIn_1(s_logisimBus2[8:0]),
.muxOut(s_logisimBus15[8:0]),
.sel(s_logisimNet3));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_5
(.carryIn(s_logisimNet16),
.carryOut(),
.dataA(s_logisimBus14[8:0]),
.dataB(s_logisimBus2[8:0]),
.result(s_logisimBus5[8:0]));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_6
(.carryIn(s_logisimNet17),
.carryOut(),
.dataA(s_logisimBus5[8:0]),
.dataB(s_logisimBus0[8:0]),
.result(s_logisimBus8[8:0]));
Comparator
#(.nrOfBits(32),
.twosComplement(1))
ARITH_7
(.aEqualsB(s_logisimNet13),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus11[31:0]),
.dataB(s_logisimBus9[31:0]));
endmodule