/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
CU
**
**
**
*****************************************************************************/
module
CU(
ALUSrc,
AlUOp,
Branch,
Jump,
MemRead,
MemWrite,
MemtoReg,
RegDst,
RegWrite,
func,
isDiv,
isMfhi,
isMflo,
isSll_shmt,
isSlti,
op_code
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[5:0]
func;
input
[5:0]
op_code;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
ALUSrc;
output
[3:0]
AlUOp;
output
Branch;
output
Jump;
output
MemRead;
output
MemWrite;
output
MemtoReg;
output
RegDst;
output
RegWrite;
output
isDiv;
output
isMfhi;
output
isMflo;
output
isSll_shmt;
output
isSlti;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[3:0]
s_logisimBus51;
wire
[5:0]
s_logisimBus52;
wire
[5:0]
s_logisimBus53;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet10;
wire
s_logisimNet11;
wire
s_logisimNet12;
wire
s_logisimNet13;
wire
s_logisimNet14;
wire
s_logisimNet15;
wire
s_logisimNet16;
wire
s_logisimNet17;
wire
s_logisimNet18;
wire
s_logisimNet19;
wire
s_logisimNet2;
wire
s_logisimNet20;
wire
s_logisimNet21;
wire
s_logisimNet22;
wire
s_logisimNet23;
wire
s_logisimNet24;
wire
s_logisimNet25;
wire
s_logisimNet26;
wire
s_logisimNet27;
wire
s_logisimNet28;
wire
s_logisimNet29;
wire
s_logisimNet3;
wire
s_logisimNet30;
wire
s_logisimNet31;
wire
s_logisimNet32;
wire
s_logisimNet33;
wire
s_logisimNet34;
wire
s_logisimNet35;
wire
s_logisimNet36;
wire
s_logisimNet37;
wire
s_logisimNet38;
wire
s_logisimNet39;
wire
s_logisimNet4;
wire
s_logisimNet40;
wire
s_logisimNet41;
wire
s_logisimNet42;
wire
s_logisimNet43;
wire
s_logisimNet44;
wire
s_logisimNet45;
wire
s_logisimNet46;
wire
s_logisimNet47;
wire
s_logisimNet48;
wire
s_logisimNet49;
wire
s_logisimNet5;
wire
s_logisimNet50;
wire
s_logisimNet6;
wire
s_logisimNet7;
wire
s_logisimNet8;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus52[5:0]
=
func;
assign
s_logisimBus53[5:0]
=
op_code;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
ALUSrc
=
s_logisimNet28;
assign
AlUOp
=
s_logisimBus51[3:0];
assign
Branch
=
s_logisimNet35;
assign
Jump
=
s_logisimNet33;
assign
MemRead
=
s_logisimNet26;
assign
MemWrite
=
s_logisimNet27;
assign
MemtoReg
=
s_logisimNet26;
assign
RegDst
=
s_logisimNet1;
assign
RegWrite
=
s_logisimNet7;
assign
isDiv
=
s_logisimNet36;
assign
isMfhi
=
s_logisimNet4;
assign
isMflo
=
s_logisimNet37;
assign
isSll_shmt
=
s_logisimNet41;
assign
isSlti
=
s_logisimNet43;
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimNet30
=
~s_logisimNet36;
assign
s_logisimNet19
=
~s_logisimBus52[5];
assign
s_logisimNet8
=
~s_logisimBus52[4];
assign
s_logisimNet16
=
~s_logisimBus52[3];
assign
s_logisimNet6
=
~s_logisimBus52[2];
assign
s_logisimNet25
=
~s_logisimBus52[1];
assign
s_logisimNet9
=
~s_logisimBus52[0];
assign
s_logisimNet24
=
~s_logisimBus53[5];
assign
s_logisimNet13
=
~s_logisimBus53[4];
assign
s_logisimNet31
=
~s_logisimBus53[3];
assign
s_logisimNet18
=
~s_logisimBus53[2];
assign
s_logisimNet10
=
~s_logisimBus53[1];
assign
s_logisimNet0
=
~s_logisimBus53[0];
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE_5_INPUTS
#(.BubblesMask({1'b0,
4'h0}))
GATES_1
(.input1(s_logisimNet27),
.input2(s_logisimNet23),
.input3(1'b0),
.input4(s_logisimNet26),
.input5(s_logisimNet43),
.result(s_logisimNet28));
OR_GATE_5_INPUTS
#(.BubblesMask({1'b0,
4'h0}))
GATES_2
(.input1(s_logisimNet1),
.input2(s_logisimNet26),
.input3(1'b0),
.input4(s_logisimNet23),
.input5(s_logisimNet43),
.result(s_logisimNet44));
AND_GATE
#(.BubblesMask(2'b00))
GATES_3
(.input1(s_logisimNet44),
.input2(s_logisimNet30),
.result(s_logisimNet7));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
mfloo
(.input1(s_logisimNet1),
.input2(s_logisimNet9),
.input3(s_logisimBus52[1]),
.input4(s_logisimNet6),
.input5(s_logisimNet16),
.input6(s_logisimBus52[4]),
.input7(s_logisimNet19),
.result(s_logisimNet37));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
div
(.input1(s_logisimNet1),
.input2(s_logisimNet9),
.input3(s_logisimBus52[1]),
.input4(s_logisimNet6),
.input5(s_logisimBus52[3]),
.input6(s_logisimBus52[4]),
.input7(s_logisimNet19),
.result(s_logisimNet36));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
sll_old
(.input1(s_logisimNet1),
.input2(s_logisimNet9),
.input3(s_logisimNet25),
.input4(s_logisimBus52[2]),
.input5(s_logisimNet16),
.input6(s_logisimNet8),
.input7(s_logisimNet19),
.result(s_logisimNet48));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
add
(.input1(s_logisimNet1),
.input2(s_logisimNet9),
.input3(s_logisimNet25),
.input4(s_logisimNet6),
.input5(s_logisimNet16),
.input6(s_logisimNet8),
.input7(s_logisimBus52[5]),
.result(s_logisimNet42));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
sub
(.input1(s_logisimNet1),
.input2(s_logisimNet9),
.input3(s_logisimBus52[1]),
.input4(s_logisimNet6),
.input5(s_logisimNet16),
.input6(s_logisimNet8),
.input7(s_logisimBus52[5]),
.result(s_logisimNet17));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
annd
(.input1(s_logisimNet1),
.input2(s_logisimNet9),
.input3(s_logisimNet25),
.input4(s_logisimBus52[2]),
.input5(s_logisimNet16),
.input6(s_logisimNet8),
.input7(s_logisimBus52[5]),
.result(s_logisimNet32));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
Or1
(.input1(s_logisimNet1),
.input2(s_logisimBus52[0]),
.input3(s_logisimNet25),
.input4(s_logisimBus52[2]),
.input5(s_logisimNet16),
.input6(s_logisimNet8),
.input7(s_logisimBus52[5]),
.result(s_logisimNet46));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
xor1
(.input1(s_logisimNet1),
.input2(s_logisimNet9),
.input3(s_logisimBus52[1]),
.input4(s_logisimBus52[2]),
.input5(s_logisimNet16),
.input6(s_logisimNet8),
.input7(s_logisimBus52[5]),
.result(s_logisimNet39));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
sll_SH
(.input1(s_logisimNet1),
.input2(s_logisimNet9),
.input3(s_logisimNet25),
.input4(s_logisimNet6),
.input5(s_logisimNet16),
.input6(s_logisimNet8),
.input7(s_logisimNet19),
.result(s_logisimNet41));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
srl1
(.input1(s_logisimNet1),
.input2(s_logisimNet9),
.input3(s_logisimBus52[1]),
.input4(s_logisimBus52[2]),
.input5(s_logisimNet16),
.input6(s_logisimNet8),
.input7(s_logisimNet19),
.result(s_logisimNet38));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
sra1
(.input1(s_logisimNet1),
.input2(s_logisimBus52[0]),
.input3(s_logisimBus52[1]),
.input4(s_logisimBus52[2]),
.input5(s_logisimNet16),
.input6(s_logisimNet8),
.input7(s_logisimNet19),
.result(s_logisimNet49));
AND_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
mfhii
(.input1(s_logisimNet1),
.input2(s_logisimNet9),
.input3(s_logisimNet25),
.input4(s_logisimNet6),
.input5(s_logisimNet16),
.input6(s_logisimBus52[4]),
.input7(s_logisimNet19),
.result(s_logisimNet4));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
R_type
(.input1(s_logisimNet0),
.input2(s_logisimNet10),
.input3(s_logisimNet18),
.input4(s_logisimNet31),
.input5(s_logisimNet13),
.input6(s_logisimNet24),
.result(s_logisimNet1));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
addi
(.input1(s_logisimNet0),
.input2(s_logisimNet10),
.input3(s_logisimNet18),
.input4(s_logisimBus53[3]),
.input5(s_logisimNet13),
.input6(s_logisimNet24),
.result(s_logisimNet23));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
sw
(.input1(s_logisimBus53[0]),
.input2(s_logisimBus53[1]),
.input3(s_logisimNet18),
.input4(s_logisimBus53[3]),
.input5(s_logisimNet13),
.input6(s_logisimBus53[5]),
.result(s_logisimNet27));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
lw
(.input1(s_logisimBus53[5]),
.input2(s_logisimNet13),
.input3(s_logisimNet31),
.input4(s_logisimNet18),
.input5(s_logisimBus53[1]),
.input6(s_logisimBus53[0]),
.result(s_logisimNet26));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
bne
(.input1(s_logisimNet24),
.input2(s_logisimNet13),
.input3(s_logisimNet31),
.input4(s_logisimBus53[2]),
.input5(s_logisimNet10),
.input6(s_logisimBus53[0]),
.result(s_logisimNet35));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
slti
(.input1(s_logisimNet24),
.input2(s_logisimNet13),
.input3(s_logisimBus53[3]),
.input4(s_logisimNet18),
.input5(s_logisimBus53[1]),
.input6(s_logisimNet0),
.result(s_logisimNet43));
AND_GATE_6_INPUTS
#(.BubblesMask({2'b00,
4'h0}))
j
(.input1(s_logisimNet24),
.input2(s_logisimNet13),
.input3(s_logisimNet31),
.input4(s_logisimNet18),
.input5(s_logisimBus53[1]),
.input6(s_logisimNet0),
.result(s_logisimNet33));
OR_GATE_4_INPUTS
#(.BubblesMask(4'h0))
GATES_23
(.input1(s_logisimNet38),
.input2(s_logisimNet49),
.input3(s_logisimNet36),
.input4(s_logisimNet39),
.result(s_logisimBus51[1]));
OR_GATE_3_INPUTS
#(.BubblesMask(3'b000))
GATES_24
(.input1(s_logisimNet32),
.input2(s_logisimNet46),
.input3(s_logisimNet39),
.result(s_logisimBus51[2]));
OR_GATE_4_INPUTS
#(.BubblesMask(4'h0))
GATES_25
(.input1(s_logisimNet48),
.input2(s_logisimNet49),
.input3(s_logisimNet38),
.input4(s_logisimNet41),
.result(s_logisimBus51[3]));
OR_GATE_8_INPUTS
#(.BubblesMask(8'h00))
GATES_26
(.input1(s_logisimNet46),
.input2(s_logisimNet35),
.input3(s_logisimNet36),
.input4(s_logisimNet17),
.input5(s_logisimNet41),
.input6(s_logisimNet49),
.input7(s_logisimNet48),
.input8(s_logisimNet43),
.result(s_logisimBus51[0]));
endmodule