/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
main
**
**
**
*****************************************************************************/
module
main(
InstDone,
Jen,
Jin,
Jout,
R1,
R10,
R11,
R12,
R13,
R14,
R15,
R16,
R17,
R18,
R19,
R2,
R20,
R21,
R22,
R23,
R24,
R25,
R26,
R27,
R28,
R29,
R3,
R30,
R31,
R4,
R5,
R6,
R7,
R8,
R9,
clk,
rst
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
Jen;
input
[31:0]
Jin;
input
clk;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
InstDone;
output
[31:0]
Jout;
output
[31:0]
R1;
output
[31:0]
R10;
output
[31:0]
R11;
output
[31:0]
R12;
output
[31:0]
R13;
output
[31:0]
R14;
output
[31:0]
R15;
output
[31:0]
R16;
output
[31:0]
R17;
output
[31:0]
R18;
output
[31:0]
R19;
output
[31:0]
R2;
output
[31:0]
R20;
output
[31:0]
R21;
output
[31:0]
R22;
output
[31:0]
R23;
output
[31:0]
R24;
output
[31:0]
R25;
output
[31:0]
R26;
output
[31:0]
R27;
output
[31:0]
R28;
output
[31:0]
R29;
output
[31:0]
R3;
output
[31:0]
R30;
output
[31:0]
R31;
output
[31:0]
R4;
output
[31:0]
R5;
output
[31:0]
R6;
output
[31:0]
R7;
output
[31:0]
R8;
output
[31:0]
R9;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus1;
wire
[31:0]
s_logisimBus10;
wire
[31:0]
s_logisimBus11;
wire
[31:0]
s_logisimBus12;
wire
[31:0]
s_logisimBus13;
wire
[31:0]
s_logisimBus14;
wire
[31:0]
s_logisimBus15;
wire
[31:0]
s_logisimBus16;
wire
[31:0]
s_logisimBus17;
wire
[31:0]
s_logisimBus18;
wire
[31:0]
s_logisimBus19;
wire
[31:0]
s_logisimBus2;
wire
[4:0]
s_logisimBus20;
wire
[4:0]
s_logisimBus21;
wire
[8:0]
s_logisimBus22;
wire
[31:0]
s_logisimBus25;
wire
[31:0]
s_logisimBus27;
wire
[31:0]
s_logisimBus29;
wire
[31:0]
s_logisimBus3;
wire
[5:0]
s_logisimBus32;
wire
[31:0]
s_logisimBus33;
wire
[31:0]
s_logisimBus34;
wire
[31:0]
s_logisimBus37;
wire
[31:0]
s_logisimBus38;
wire
[31:0]
s_logisimBus4;
wire
[31:0]
s_logisimBus40;
wire
[31:0]
s_logisimBus42;
wire
[31:0]
s_logisimBus43;
wire
[31:0]
s_logisimBus44;
wire
[31:0]
s_logisimBus45;
wire
[31:0]
s_logisimBus46;
wire
[31:0]
s_logisimBus47;
wire
[31:0]
s_logisimBus48;
wire
[31:0]
s_logisimBus49;
wire
[31:0]
s_logisimBus5;
wire
[31:0]
s_logisimBus50;
wire
[31:0]
s_logisimBus51;
wire
[31:0]
s_logisimBus52;
wire
[31:0]
s_logisimBus53;
wire
[31:0]
s_logisimBus54;
wire
[31:0]
s_logisimBus55;
wire
[31:0]
s_logisimBus56;
wire
[31:0]
s_logisimBus57;
wire
[31:0]
s_logisimBus58;
wire
[4:0]
s_logisimBus59;
wire
[31:0]
s_logisimBus6;
wire
[4:0]
s_logisimBus60;
wire
[31:0]
s_logisimBus61;
wire
[31:0]
s_logisimBus65;
wire
[8:0]
s_logisimBus68;
wire
[31:0]
s_logisimBus69;
wire
[31:0]
s_logisimBus7;
wire
[31:0]
s_logisimBus71;
wire
[31:0]
s_logisimBus73;
wire
[31:0]
s_logisimBus76;
wire
[31:0]
s_logisimBus8;
wire
[4:0]
s_logisimBus82;
wire
[4:0]
s_logisimBus83;
wire
[31:0]
s_logisimBus84;
wire
[31:0]
s_logisimBus85;
wire
[3:0]
s_logisimBus86;
wire
[5:0]
s_logisimBus87;
wire
[4:0]
s_logisimBus88;
wire
[31:0]
s_logisimBus9;
wire
[15:0]
s_logisimBus91;
wire
s_logisimNet23;
wire
s_logisimNet24;
wire
s_logisimNet26;
wire
s_logisimNet28;
wire
s_logisimNet30;
wire
s_logisimNet31;
wire
s_logisimNet35;
wire
s_logisimNet36;
wire
s_logisimNet41;
wire
s_logisimNet62;
wire
s_logisimNet63;
wire
s_logisimNet64;
wire
s_logisimNet66;
wire
s_logisimNet67;
wire
s_logisimNet70;
wire
s_logisimNet72;
wire
s_logisimNet74;
wire
s_logisimNet75;
wire
s_logisimNet77;
wire
s_logisimNet78;
wire
s_logisimNet79;
wire
s_logisimNet80;
wire
s_logisimNet81;
wire
s_logisimNet89;
wire
s_logisimNet90;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus1[31:0]
=
Jin;
assign
s_logisimNet31
=
Jen;
assign
s_logisimNet81
=
rst;
assign
s_logisimNet89
=
clk;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
InstDone
=
s_logisimNet64;
assign
Jout
=
s_logisimBus3[31:0];
assign
R1
=
s_logisimBus45[31:0];
assign
R10
=
s_logisimBus8[31:0];
assign
R11
=
s_logisimBus48[31:0];
assign
R12
=
s_logisimBus9[31:0];
assign
R13
=
s_logisimBus49[31:0];
assign
R14
=
s_logisimBus10[31:0];
assign
R15
=
s_logisimBus50[31:0];
assign
R16
=
s_logisimBus11[31:0];
assign
R17
=
s_logisimBus51[31:0];
assign
R18
=
s_logisimBus12[31:0];
assign
R19
=
s_logisimBus52[31:0];
assign
R2
=
s_logisimBus6[31:0];
assign
R20
=
s_logisimBus13[31:0];
assign
R21
=
s_logisimBus53[31:0];
assign
R22
=
s_logisimBus14[31:0];
assign
R23
=
s_logisimBus54[31:0];
assign
R24
=
s_logisimBus15[31:0];
assign
R25
=
s_logisimBus55[31:0];
assign
R26
=
s_logisimBus16[31:0];
assign
R27
=
s_logisimBus56[31:0];
assign
R28
=
s_logisimBus17[31:0];
assign
R29
=
s_logisimBus57[31:0];
assign
R3
=
s_logisimBus44[31:0];
assign
R30
=
s_logisimBus18[31:0];
assign
R31
=
s_logisimBus58[31:0];
assign
R4
=
s_logisimBus5[31:0];
assign
R5
=
s_logisimBus46[31:0];
assign
R6
=
s_logisimBus7[31:0];
assign
R7
=
s_logisimBus43[31:0];
assign
R8
=
s_logisimBus4[31:0];
assign
R9
=
s_logisimBus47[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus76[31:0]
=
32'h00000000;
assign
s_logisimBus59[4:0]
=
{1'b0,
4'h0};
assign
s_logisimBus34[0]
=
s_logisimNet30;
assign
s_logisimBus34[1]
=
1'b0;
assign
s_logisimBus34[2]
=
1'b0;
assign
s_logisimBus34[3]
=
1'b0;
assign
s_logisimBus34[4]
=
1'b0;
assign
s_logisimBus34[5]
=
1'b0;
assign
s_logisimBus34[6]
=
1'b0;
assign
s_logisimBus34[7]
=
1'b0;
assign
s_logisimBus34[8]
=
1'b0;
assign
s_logisimBus34[9]
=
1'b0;
assign
s_logisimBus34[10]
=
1'b0;
assign
s_logisimBus34[11]
=
1'b0;
assign
s_logisimBus34[12]
=
1'b0;
assign
s_logisimBus34[13]
=
1'b0;
assign
s_logisimBus34[14]
=
1'b0;
assign
s_logisimBus34[15]
=
1'b0;
assign
s_logisimBus34[16]
=
1'b0;
assign
s_logisimBus34[17]
=
1'b0;
assign
s_logisimBus34[18]
=
1'b0;
assign
s_logisimBus34[19]
=
1'b0;
assign
s_logisimBus34[20]
=
1'b0;
assign
s_logisimBus34[21]
=
1'b0;
assign
s_logisimBus34[22]
=
1'b0;
assign
s_logisimBus34[23]
=
1'b0;
assign
s_logisimBus34[24]
=
1'b0;
assign
s_logisimBus34[25]
=
1'b0;
assign
s_logisimBus34[26]
=
1'b0;
assign
s_logisimBus34[27]
=
1'b0;
assign
s_logisimBus34[28]
=
1'b0;
assign
s_logisimBus34[29]
=
1'b0;
assign
s_logisimBus34[30]
=
1'b0;
assign
s_logisimBus34[31]
=
1'b0;
assign
s_logisimNet77
=
1'b1;
assign
s_logisimBus69[0]
=
s_logisimBus91[0];
assign
s_logisimBus69[1]
=
s_logisimBus91[1];
assign
s_logisimBus69[2]
=
s_logisimBus91[2];
assign
s_logisimBus69[3]
=
s_logisimBus91[3];
assign
s_logisimBus69[4]
=
s_logisimBus91[4];
assign
s_logisimBus69[5]
=
s_logisimBus91[5];
assign
s_logisimBus69[6]
=
s_logisimBus91[6];
assign
s_logisimBus69[7]
=
s_logisimBus91[7];
assign
s_logisimBus69[8]
=
s_logisimBus91[8];
assign
s_logisimBus69[9]
=
s_logisimBus91[9];
assign
s_logisimBus69[10]
=
s_logisimBus91[10];
assign
s_logisimBus69[11]
=
s_logisimBus91[11];
assign
s_logisimBus69[12]
=
s_logisimBus91[12];
assign
s_logisimBus69[13]
=
s_logisimBus91[13];
assign
s_logisimBus69[14]
=
s_logisimBus91[14];
assign
s_logisimBus69[15]
=
s_logisimBus91[15];
assign
s_logisimBus69[16]
=
s_logisimBus91[15];
assign
s_logisimBus69[17]
=
s_logisimBus91[15];
assign
s_logisimBus69[18]
=
s_logisimBus91[15];
assign
s_logisimBus69[19]
=
s_logisimBus91[15];
assign
s_logisimBus69[20]
=
s_logisimBus91[15];
assign
s_logisimBus69[21]
=
s_logisimBus91[15];
assign
s_logisimBus69[22]
=
s_logisimBus91[15];
assign
s_logisimBus69[23]
=
s_logisimBus91[15];
assign
s_logisimBus69[24]
=
s_logisimBus91[15];
assign
s_logisimBus69[25]
=
s_logisimBus91[15];
assign
s_logisimBus69[26]
=
s_logisimBus91[15];
assign
s_logisimBus69[27]
=
s_logisimBus91[15];
assign
s_logisimBus69[28]
=
s_logisimBus91[15];
assign
s_logisimBus69[29]
=
s_logisimBus91[15];
assign
s_logisimBus69[30]
=
s_logisimBus91[15];
assign
s_logisimBus69[31]
=
s_logisimBus91[15];
assign
s_logisimBus61[0]
=
s_logisimBus21[0];
assign
s_logisimBus61[1]
=
s_logisimBus21[1];
assign
s_logisimBus61[2]
=
s_logisimBus21[2];
assign
s_logisimBus61[3]
=
s_logisimBus21[3];
assign
s_logisimBus61[4]
=
s_logisimBus21[4];
assign
s_logisimBus61[5]
=
s_logisimBus21[4];
assign
s_logisimBus61[6]
=
s_logisimBus21[4];
assign
s_logisimBus61[7]
=
s_logisimBus21[4];
assign
s_logisimBus61[8]
=
s_logisimBus21[4];
assign
s_logisimBus61[9]
=
s_logisimBus21[4];
assign
s_logisimBus61[10]
=
s_logisimBus21[4];
assign
s_logisimBus61[11]
=
s_logisimBus21[4];
assign
s_logisimBus61[12]
=
s_logisimBus21[4];
assign
s_logisimBus61[13]
=
s_logisimBus21[4];
assign
s_logisimBus61[14]
=
s_logisimBus21[4];
assign
s_logisimBus61[15]
=
s_logisimBus21[4];
assign
s_logisimBus61[16]
=
s_logisimBus21[4];
assign
s_logisimBus61[17]
=
s_logisimBus21[4];
assign
s_logisimBus61[18]
=
s_logisimBus21[4];
assign
s_logisimBus61[19]
=
s_logisimBus21[4];
assign
s_logisimBus61[20]
=
s_logisimBus21[4];
assign
s_logisimBus61[21]
=
s_logisimBus21[4];
assign
s_logisimBus61[22]
=
s_logisimBus21[4];
assign
s_logisimBus61[23]
=
s_logisimBus21[4];
assign
s_logisimBus61[24]
=
s_logisimBus21[4];
assign
s_logisimBus61[25]
=
s_logisimBus21[4];
assign
s_logisimBus61[26]
=
s_logisimBus21[4];
assign
s_logisimBus61[27]
=
s_logisimBus21[4];
assign
s_logisimBus61[28]
=
s_logisimBus21[4];
assign
s_logisimBus61[29]
=
s_logisimBus21[4];
assign
s_logisimBus61[30]
=
s_logisimBus21[4];
assign
s_logisimBus61[31]
=
s_logisimBus21[4];
assign
s_logisimNet79
=
1'b0;
assign
s_logisimNet80
=
1'b0;
assign
s_logisimNet64
=
~s_logisimNet28;
assign
s_logisimNet72
=
~s_logisimNet62;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE
#(.BubblesMask(2'b00))
GATES_1
(.input1(s_logisimNet72),
.input2(s_logisimNet63),
.result(s_logisimNet28));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus83[4:0]),
.muxIn_1(s_logisimBus88[4:0]),
.muxOut(s_logisimBus20[4:0]),
.sel(s_logisimNet35));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus59[4:0]),
.muxIn_1(s_logisimBus20[4:0]),
.muxOut(s_logisimBus60[4:0]),
.sel(s_logisimNet74));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus71[31:0]),
.muxIn_1(s_logisimBus27[31:0]),
.muxOut(s_logisimBus0[31:0]),
.sel(s_logisimNet67));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus0[31:0]),
.muxIn_1(s_logisimBus34[31:0]),
.muxOut(s_logisimBus65[31:0]),
.sel(s_logisimNet41));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus65[31:0]),
.muxIn_1(s_logisimBus73[31:0]),
.muxOut(s_logisimBus2[31:0]),
.sel(s_logisimNet66));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_7
(.enable(1'b1),
.muxIn_0(s_logisimBus2[31:0]),
.muxIn_1(s_logisimBus42[31:0]),
.muxOut(s_logisimBus38[31:0]),
.sel(s_logisimNet75));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus85[31:0]),
.muxIn_1(s_logisimBus69[31:0]),
.muxOut(s_logisimBus37[31:0]),
.sel(s_logisimNet23));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_9
(.enable(1'b1),
.muxIn_0(s_logisimBus37[31:0]),
.muxIn_1(s_logisimBus61[31:0]),
.muxOut(s_logisimBus40[31:0]),
.sel(s_logisimNet26));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_10
(.enable(1'b1),
.muxIn_0(s_logisimBus84[31:0]),
.muxIn_1(s_logisimBus85[31:0]),
.muxOut(s_logisimBus19[31:0]),
.sel(s_logisimNet26));
Comparator
#(.nrOfBits(32),
.twosComplement(1))
ARITH_11
(.aEqualsB(),
.aGreaterThanB(s_logisimNet30),
.aLessThanB(),
.dataA(s_logisimBus76[31:0]),
.dataB(s_logisimBus71[31:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
programCounter
(.clock(s_logisimNet89),
.clockEnable(s_logisimNet77),
.d(s_logisimBus22[8:0]),
.q(s_logisimBus68[8:0]),
.reset(s_logisimNet81),
.tick(1'b1));
D_FLIPFLOP
#(.invertClockEnable(0))
MEMORY_13
(.clock(s_logisimNet89),
.d(s_logisimNet78),
.preset(1'b0),
.q(s_logisimNet62),
.qBar(),
.reset(s_logisimNet81),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_14
(.clock(s_logisimNet89),
.clockEnable(s_logisimNet63),
.d(s_logisimBus71[31:0]),
.q(s_logisimBus73[31:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_15
(.clock(s_logisimNet89),
.clockEnable(s_logisimNet63),
.d(s_logisimBus33[31:0]),
.q(s_logisimBus42[31:0]),
.reset(1'b0),
.tick(1'b1));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
ALU
ALU_1
(.a(s_logisimBus19[31:0]),
.aluop(s_logisimBus86[3:0]),
.b(s_logisimBus40[31:0]),
.clk(s_logisimNet89),
.done(s_logisimNet78),
.output_inc(s_logisimNet79),
.output_inverted(s_logisimNet80),
.res_high(s_logisimBus33[31:0]),
.res_low(s_logisimBus71[31:0]),
.rst(s_logisimNet81));
regfile
RF
(.Aread0(s_logisimBus82[4:0]),
.Aread1(s_logisimBus83[4:0]),
.Awrite(s_logisimBus60[4:0]),
.Dread0(s_logisimBus84[31:0]),
.Dread1(s_logisimBus85[31:0]),
.Dwrite(s_logisimBus38[31:0]),
.R1(s_logisimBus45[31:0]),
.R10(s_logisimBus8[31:0]),
.R11(s_logisimBus48[31:0]),
.R12(s_logisimBus9[31:0]),
.R13(s_logisimBus49[31:0]),
.R14(s_logisimBus10[31:0]),
.R15(s_logisimBus50[31:0]),
.R16(s_logisimBus11[31:0]),
.R17(s_logisimBus51[31:0]),
.R18(s_logisimBus12[31:0]),
.R19(s_logisimBus52[31:0]),
.R2(s_logisimBus6[31:0]),
.R20(s_logisimBus13[31:0]),
.R21(s_logisimBus53[31:0]),
.R22(s_logisimBus14[31:0]),
.R23(s_logisimBus54[31:0]),
.R24(s_logisimBus15[31:0]),
.R25(s_logisimBus55[31:0]),
.R26(s_logisimBus16[31:0]),
.R27(s_logisimBus56[31:0]),
.R28(s_logisimBus17[31:0]),
.R29(s_logisimBus57[31:0]),
.R3(s_logisimBus44[31:0]),
.R30(s_logisimBus18[31:0]),
.R31(s_logisimBus58[31:0]),
.R4(s_logisimBus5[31:0]),
.R5(s_logisimBus46[31:0]),
.R6(s_logisimBus7[31:0]),
.R7(s_logisimBus43[31:0]),
.R8(s_logisimBus4[31:0]),
.R9(s_logisimBus47[31:0]),
.clk(s_logisimNet89),
.rst(s_logisimNet81));
CU
Control_Unit
(.ALUSrc(s_logisimNet23),
.AlUOp(s_logisimBus86[3:0]),
.Branch(s_logisimNet90),
.Jump(s_logisimNet70),
.MemRead(s_logisimNet24),
.MemWrite(s_logisimNet36),
.MemtoReg(s_logisimNet67),
.RegDst(s_logisimNet35),
.RegWrite(s_logisimNet74),
.func(s_logisimBus87[5:0]),
.isDiv(s_logisimNet63),
.isMfhi(s_logisimNet75),
.isMflo(s_logisimNet66),
.isSll_shmt(s_logisimNet26),
.isSlti(s_logisimNet41),
.op_code(s_logisimBus32[5:0]));
INC_decoder
INC
(.fuunc(s_logisimBus87[5:0]),
.imm(s_logisimBus91[15:0]),
.inc(s_logisimBus29[31:0]),
.op(s_logisimBus32[5:0]),
.rd(s_logisimBus88[4:0]),
.rs(s_logisimBus82[4:0]),
.rt(s_logisimBus83[4:0]),
.shamt(s_logisimBus21[4:0]));
jtag_ram512
I_mem
(.Addr(s_logisimBus68[8:0]),
.Din(32'd0),
.Dout(s_logisimBus29[31:0]),
.Jen(s_logisimNet31),
.Jin(s_logisimBus1[31:0]),
.Jout(s_logisimBus25[31:0]),
.Wen(1'b0),
.clk(s_logisimNet89));
jtag_ram512
D_mem
(.Addr(s_logisimBus71[8:0]),
.Din(s_logisimBus85[31:0]),
.Dout(s_logisimBus27[31:0]),
.Jen(s_logisimNet31),
.Jin(s_logisimBus25[31:0]),
.Jout(s_logisimBus3[31:0]),
.Wen(s_logisimNet36),
.clk(s_logisimNet89));
PC_Update
PC_Update_1
(.Branch(s_logisimNet90),
.Eq(s_logisimBus71[31:0]),
.Imm(s_logisimBus91[15:0]),
.Jump(s_logisimNet70),
.PC(s_logisimBus68[8:0]),
.PC_out(s_logisimBus22[8:0]),
.divIsActive(s_logisimNet28));
endmodule