/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
ALU
**
**
**
*****************************************************************************/
module
ALU(
a,
aluop,
b,
clk,
done,
output_inc,
output_inverted,
res_high,
res_low,
rst
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[3:0]
aluop;
input
[31:0]
b;
input
clk;
input
output_inc;
input
output_inverted;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
done;
output
[31:0]
res_high;
output
[31:0]
res_low;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus1;
wire
[63:0]
s_logisimBus11;
wire
[31:0]
s_logisimBus12;
wire
[63:0]
s_logisimBus14;
wire
[63:0]
s_logisimBus16;
wire
[63:0]
s_logisimBus18;
wire
[63:0]
s_logisimBus19;
wire
[31:0]
s_logisimBus20;
wire
[63:0]
s_logisimBus23;
wire
[63:0]
s_logisimBus24;
wire
[63:0]
s_logisimBus26;
wire
[3:0]
s_logisimBus28;
wire
[63:0]
s_logisimBus29;
wire
[31:0]
s_logisimBus30;
wire
[63:0]
s_logisimBus31;
wire
[63:0]
s_logisimBus35;
wire
[63:0]
s_logisimBus36;
wire
[63:0]
s_logisimBus37;
wire
[31:0]
s_logisimBus38;
wire
[63:0]
s_logisimBus39;
wire
[31:0]
s_logisimBus40;
wire
[63:0]
s_logisimBus41;
wire
[31:0]
s_logisimBus42;
wire
[63:0]
s_logisimBus44;
wire
[63:0]
s_logisimBus5;
wire
[63:0]
s_logisimBus9;
wire
s_logisimNet13;
wire
s_logisimNet22;
wire
s_logisimNet32;
wire
s_logisimNet33;
wire
s_logisimNet34;
wire
s_logisimNet43;
wire
s_logisimNet45;
wire
s_logisimNet7;
wire
s_logisimNet8;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
wiring
is
defined
**
*******************************************************************************/
assign
s_logisimBus16[32]
=
s_logisimBus20[0];
assign
s_logisimBus16[33]
=
s_logisimBus20[1];
assign
s_logisimBus16[34]
=
s_logisimBus20[2];
assign
s_logisimBus16[35]
=
s_logisimBus20[3];
assign
s_logisimBus16[36]
=
s_logisimBus20[4];
assign
s_logisimBus16[37]
=
s_logisimBus20[5];
assign
s_logisimBus16[38]
=
s_logisimBus20[6];
assign
s_logisimBus16[39]
=
s_logisimBus20[7];
assign
s_logisimBus16[40]
=
s_logisimBus20[8];
assign
s_logisimBus16[41]
=
s_logisimBus20[9];
assign
s_logisimBus16[42]
=
s_logisimBus20[10];
assign
s_logisimBus16[43]
=
s_logisimBus20[11];
assign
s_logisimBus16[44]
=
s_logisimBus20[12];
assign
s_logisimBus16[45]
=
s_logisimBus20[13];
assign
s_logisimBus16[46]
=
s_logisimBus20[14];
assign
s_logisimBus16[47]
=
s_logisimBus20[15];
assign
s_logisimBus16[48]
=
s_logisimBus20[16];
assign
s_logisimBus16[49]
=
s_logisimBus20[17];
assign
s_logisimBus16[50]
=
s_logisimBus20[18];
assign
s_logisimBus16[51]
=
s_logisimBus20[19];
assign
s_logisimBus16[52]
=
s_logisimBus20[20];
assign
s_logisimBus16[53]
=
s_logisimBus20[21];
assign
s_logisimBus16[54]
=
s_logisimBus20[22];
assign
s_logisimBus16[55]
=
s_logisimBus20[23];
assign
s_logisimBus16[56]
=
s_logisimBus20[24];
assign
s_logisimBus16[57]
=
s_logisimBus20[25];
assign
s_logisimBus16[58]
=
s_logisimBus20[26];
assign
s_logisimBus16[59]
=
s_logisimBus20[27];
assign
s_logisimBus16[60]
=
s_logisimBus20[28];
assign
s_logisimBus16[61]
=
s_logisimBus20[29];
assign
s_logisimBus16[62]
=
s_logisimBus20[30];
assign
s_logisimBus16[63]
=
s_logisimBus20[31];
assign
s_logisimBus29[32]
=
s_logisimBus20[0];
assign
s_logisimBus29[33]
=
s_logisimBus20[1];
assign
s_logisimBus29[34]
=
s_logisimBus20[2];
assign
s_logisimBus29[35]
=
s_logisimBus20[3];
assign
s_logisimBus29[36]
=
s_logisimBus20[4];
assign
s_logisimBus29[37]
=
s_logisimBus20[5];
assign
s_logisimBus29[38]
=
s_logisimBus20[6];
assign
s_logisimBus29[39]
=
s_logisimBus20[7];
assign
s_logisimBus29[40]
=
s_logisimBus20[8];
assign
s_logisimBus29[41]
=
s_logisimBus20[9];
assign
s_logisimBus29[42]
=
s_logisimBus20[10];
assign
s_logisimBus29[43]
=
s_logisimBus20[11];
assign
s_logisimBus29[44]
=
s_logisimBus20[12];
assign
s_logisimBus29[45]
=
s_logisimBus20[13];
assign
s_logisimBus29[46]
=
s_logisimBus20[14];
assign
s_logisimBus29[47]
=
s_logisimBus20[15];
assign
s_logisimBus29[48]
=
s_logisimBus20[16];
assign
s_logisimBus29[49]
=
s_logisimBus20[17];
assign
s_logisimBus29[50]
=
s_logisimBus20[18];
assign
s_logisimBus29[51]
=
s_logisimBus20[19];
assign
s_logisimBus29[52]
=
s_logisimBus20[20];
assign
s_logisimBus29[53]
=
s_logisimBus20[21];
assign
s_logisimBus29[54]
=
s_logisimBus20[22];
assign
s_logisimBus29[55]
=
s_logisimBus20[23];
assign
s_logisimBus29[56]
=
s_logisimBus20[24];
assign
s_logisimBus29[57]
=
s_logisimBus20[25];
assign
s_logisimBus29[58]
=
s_logisimBus20[26];
assign
s_logisimBus29[59]
=
s_logisimBus20[27];
assign
s_logisimBus29[60]
=
s_logisimBus20[28];
assign
s_logisimBus29[61]
=
s_logisimBus20[29];
assign
s_logisimBus29[62]
=
s_logisimBus20[30];
assign
s_logisimBus29[63]
=
s_logisimBus20[31];
assign
s_logisimBus41[32]
=
s_logisimBus20[0];
assign
s_logisimBus41[33]
=
s_logisimBus20[1];
assign
s_logisimBus41[34]
=
s_logisimBus20[2];
assign
s_logisimBus41[35]
=
s_logisimBus20[3];
assign
s_logisimBus41[36]
=
s_logisimBus20[4];
assign
s_logisimBus41[37]
=
s_logisimBus20[5];
assign
s_logisimBus41[38]
=
s_logisimBus20[6];
assign
s_logisimBus41[39]
=
s_logisimBus20[7];
assign
s_logisimBus41[40]
=
s_logisimBus20[8];
assign
s_logisimBus41[41]
=
s_logisimBus20[9];
assign
s_logisimBus41[42]
=
s_logisimBus20[10];
assign
s_logisimBus41[43]
=
s_logisimBus20[11];
assign
s_logisimBus41[44]
=
s_logisimBus20[12];
assign
s_logisimBus41[45]
=
s_logisimBus20[13];
assign
s_logisimBus41[46]
=
s_logisimBus20[14];
assign
s_logisimBus41[47]
=
s_logisimBus20[15];
assign
s_logisimBus41[48]
=
s_logisimBus20[16];
assign
s_logisimBus41[49]
=
s_logisimBus20[17];
assign
s_logisimBus41[50]
=
s_logisimBus20[18];
assign
s_logisimBus41[51]
=
s_logisimBus20[19];
assign
s_logisimBus41[52]
=
s_logisimBus20[20];
assign
s_logisimBus41[53]
=
s_logisimBus20[21];
assign
s_logisimBus41[54]
=
s_logisimBus20[22];
assign
s_logisimBus41[55]
=
s_logisimBus20[23];
assign
s_logisimBus41[56]
=
s_logisimBus20[24];
assign
s_logisimBus41[57]
=
s_logisimBus20[25];
assign
s_logisimBus41[58]
=
s_logisimBus20[26];
assign
s_logisimBus41[59]
=
s_logisimBus20[27];
assign
s_logisimBus41[60]
=
s_logisimBus20[28];
assign
s_logisimBus41[61]
=
s_logisimBus20[29];
assign
s_logisimBus41[62]
=
s_logisimBus20[30];
assign
s_logisimBus41[63]
=
s_logisimBus20[31];
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus28[3:0]
=
aluop;
assign
s_logisimBus38[31:0]
=
b;
assign
s_logisimBus42[31:0]
=
a;
assign
s_logisimNet32
=
output_inverted;
assign
s_logisimNet33
=
rst;
assign
s_logisimNet43
=
clk;
assign
s_logisimNet45
=
output_inc;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
done
=
s_logisimNet34;
assign
res_high
=
s_logisimBus9[63:32];
assign
res_low
=
s_logisimBus9[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimNet7
=
1'b1;
assign
s_logisimBus20[31:0]
=
32'h00000000;
assign
s_logisimNet13
=
1'b0;
assign
s_logisimBus30[31:0]
=
32'hFFFFFFFF;
assign
s_logisimBus19[63:33]
=
{3'b000,
28'h0000000};
assign
s_logisimBus12[31:0]
=
32'h00000000;
assign
s_logisimBus44[63:0]
=
64'h0000000000000000;
assign
s_logisimBus40
=
~s_logisimBus38;
assign
s_logisimBus39
=
~s_logisimBus5;
assign
s_logisimBus1
=
~s_logisimBus42;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE_BUS
#(.BubblesMask(2'b00),
.NrOfBits(32))
GATES_1
(.input1(s_logisimBus42[31:0]),
.input2(s_logisimBus38[31:0]),
.result(s_logisimBus29[31:0]));
XOR_GATE_BUS_ONEHOT
#(.BubblesMask(2'b00),
.NrOfBits(32))
GATES_2
(.input1(s_logisimBus42[31:0]),
.input2(s_logisimBus38[31:0]),
.result(s_logisimBus16[31:0]));
AND_GATE_BUS
#(.BubblesMask(2'b00),
.NrOfBits(32))
GATES_3
(.input1(s_logisimBus42[31:0]),
.input2(s_logisimBus38[31:0]),
.result(s_logisimBus41[31:0]));
Multiplexer_bus_16
#(.nrOfBits(64))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus19[63:0]),
.muxIn_1(s_logisimBus37[63:0]),
.muxIn_10(s_logisimBus23[63:0]),
.muxIn_11(s_logisimBus18[63:0]),
.muxIn_12(s_logisimBus14[63:0]),
.muxIn_13(64'd0),
.muxIn_14(64'd0),
.muxIn_15(64'd0),
.muxIn_2(s_logisimBus31[63:0]),
.muxIn_3(s_logisimBus35[63:0]),
.muxIn_4(s_logisimBus41[63:0]),
.muxIn_5(s_logisimBus29[63:0]),
.muxIn_6(s_logisimBus16[63:0]),
.muxIn_7(s_logisimBus36[63:0]),
.muxIn_8(s_logisimBus24[63:0]),
.muxIn_9(s_logisimBus26[63:0]),
.muxOut(s_logisimBus5[63:0]),
.sel(s_logisimBus28[3:0]));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus30[31:0]),
.muxIn_1(s_logisimBus12[31:0]),
.muxOut(s_logisimBus37[63:32]),
.sel(s_logisimNet8));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus5[63:0]),
.muxIn_1(s_logisimBus39[63:0]),
.muxOut(s_logisimBus11[63:0]),
.sel(s_logisimNet32));
Adder
#(.extendedBits(65),
.nrOfBits(64))
ARITH_7
(.carryIn(s_logisimNet45),
.carryOut(),
.dataA(s_logisimBus44[63:0]),
.dataB(s_logisimBus11[63:0]),
.result(s_logisimBus9[63:0]));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
ALU_MUL
ALU_MUL_1
(.a(s_logisimBus42[31:0]),
.b(s_logisimBus38[31:0]),
.mul_out(s_logisimBus31[63:0]));
ALU_CLO
ALU_CLO_1
(.A(s_logisimBus42[31:0]),
.OUTTTT(s_logisimBus36[63:0]));
ALU_CLO
ALU_CLO_2
(.A(s_logisimBus1[31:0]),
.OUTTTT(s_logisimBus24[63:0]));
ALU_DIV
ALU_DIV_1
(.clk(s_logisimNet43),
.dividend(s_logisimBus42[31:0]),
.divisor(s_logisimBus38[31:0]),
.done(s_logisimNet34),
.quotient(s_logisimBus35[31:0]),
.remainder(s_logisimBus35[63:32]));
ALU_ROTATE
ALU_ROTATE_1
(.a(s_logisimBus42[31:0]),
.b(s_logisimBus38[31:0]),
.ouuut(s_logisimBus14[63:0]));
ALU_CSA
ALU_CSA_1
(.A(s_logisimBus42[31:0]),
.B(s_logisimBus38[31:0]),
.SUM(s_logisimBus19[31:0]),
.cin(s_logisimNet13),
.cout(s_logisimBus19[32]));
ALU_CSA
ALU_CSA_2
(.A(s_logisimBus42[31:0]),
.B(s_logisimBus40[31:0]),
.SUM(s_logisimBus37[31:0]),
.cin(s_logisimNet7),
.cout(s_logisimNet8));
ALU_SRA
ALU_SRA_1
(.a(s_logisimBus42[31:0]),
.b(s_logisimBus38[31:0]),
.output1(s_logisimBus18[63:0]));
ALU_SRL
ALU_SRL_1
(.a(s_logisimBus42[31:0]),
.b(s_logisimBus38[31:0]),
.output1(s_logisimBus23[63:0]));
ALU_SLL
ALU_SLL_1
(.a(s_logisimBus42[31:0]),
.b(s_logisimBus38[31:0]),
.output1(s_logisimBus26[63:0]));
endmodule